              fgallag0x00003_0 = 
          (!fgallag_sel[2]) ? 
                       fgallag0x00002_0_q: 
                       fgallag0x00002_1_q;
              fgallag0x00003_1 = 
          (!fgallag_sel[2]) ? 
                       fgallag0x00002_2_q: 
                       fgallag0x00002_3_q;
              fgallag0x00003_2 = 
          (!fgallag_sel[2]) ? 
                       fgallag0x00002_4_q: 
                       fgallag0x00002_5_q;
              fgallag0x00003_3 = 
          (!fgallag_sel[2]) ? 
                       fgallag0x00002_6_q: 
                       fgallag0x00002_7_q;
              fgallag0x00003_4 = 
          (!fgallag_sel[2]) ? 
                       fgallag0x00002_8_q: 
                       fgallag0x00002_9_q;
              fgallag0x00003_5 = 
          (!fgallag_sel[2]) ? 
                       fgallag0x00002_10_q: 
                       fgallag0x00002_11_q;
              fgallag0x00003_6 = 
          (!fgallag_sel[2]) ? 
                       fgallag0x00002_12_q: 
                       fgallag0x00002_13_q;
              fgallag0x00003_7 = 
          (!fgallag_sel[2]) ? 
                       fgallag0x00002_14_q: 
                       fgallag0x00002_15_q;
              fgallag0x00003_8 = 
          (!fgallag_sel[2]) ? 
                       fgallag0x00002_16_q: 
                       fgallag0x00002_17_q;
              fgallag0x00003_9 = 
          (!fgallag_sel[2]) ? 
                       fgallag0x00002_18_q: 
                       fgallag0x00002_19_q;
              fgallag0x00003_10 = 
          (!fgallag_sel[2]) ? 
                       fgallag0x00002_20_q: 
                       fgallag0x00002_21_q;
              fgallag0x00003_11 = 
          (!fgallag_sel[2]) ? 
                       fgallag0x00002_22_q: 
                       fgallag0x00002_23_q;
              fgallag0x00003_12 = 
          (!fgallag_sel[2]) ? 
                       fgallag0x00002_24_q: 
                       fgallag0x00002_25_q;
              fgallag0x00003_13 = 
          (!fgallag_sel[2]) ? 
                       fgallag0x00002_26_q: 
                       fgallag0x00002_27_q;
              fgallag0x00003_14 = 
          (!fgallag_sel[2]) ? 
                       fgallag0x00002_28_q: 
                       fgallag0x00002_29_q;
              fgallag0x00003_15 = 
          (!fgallag_sel[2]) ? 
                       fgallag0x00002_30_q: 
                       fgallag0x00002_31_q;
              fgallag0x00003_16 = 
          (!fgallag_sel[2]) ? 
                       fgallag0x00002_32_q: 
                       fgallag0x00002_33_q;
              fgallag0x00003_17 = 
          (!fgallag_sel[2]) ? 
                       fgallag0x00002_34_q: 
                       fgallag0x00002_35_q;
              fgallag0x00003_18 = 
          (!fgallag_sel[2]) ? 
                       fgallag0x00002_36_q: 
                       fgallag0x00002_37_q;
              fgallag0x00003_19 = 
          (!fgallag_sel[2]) ? 
                       fgallag0x00002_38_q: 
                       fgallag0x00002_39_q;
              fgallag0x00003_20 = 
          (!fgallag_sel[2]) ? 
                       fgallag0x00002_40_q: 
                       fgallag0x00002_41_q;
              fgallag0x00003_21 = 
          (!fgallag_sel[2]) ? 
                       fgallag0x00002_42_q: 
                       fgallag0x00002_43_q;
              fgallag0x00003_22 = 
          (!fgallag_sel[2]) ? 
                       fgallag0x00002_44_q: 
                       fgallag0x00002_45_q;
               fgallag0x00003_23 =  fgallag0x00002_46_q ;
               fgallag0x00003_24 =  fgallag0x00002_48_q ;
              fgallag0x00003_25 = 
          (!fgallag_sel[2]) ? 
                       fgallag0x00002_50_q: 
                       fgallag0x00002_51_q;
              fgallag0x00003_26 = 
          (!fgallag_sel[2]) ? 
                       fgallag0x00002_52_q: 
                       fgallag0x00002_53_q;
               fgallag0x00003_27 =  fgallag0x00002_54_q ;
              fgallag0x00003_28 = 
          (!fgallag_sel[2]) ? 
                       fgallag0x00002_56_q: 
                       fgallag0x00002_57_q;
               fgallag0x00003_29 =  fgallag0x00002_58_q ;
               fgallag0x00003_30 =  fgallag0x00002_60_q ;
              fgallag0x00003_31 = 
          (!fgallag_sel[2]) ? 
                       fgallag0x00002_62_q: 
                       fgallag0x00002_63_q;
               fgallag0x00003_32 =  fgallag0x00002_64_q ;
               fgallag0x00003_33 =  fgallag0x00002_66_q ;
               fgallag0x00003_34 =  fgallag0x00002_68_q ;
              fgallag0x00003_35 = 
          (!fgallag_sel[2]) ? 
                       fgallag0x00002_70_q: 
                       fgallag0x00002_71_q;
               fgallag0x00003_36 =  fgallag0x00002_72_q ;
               fgallag0x00003_37 =  fgallag0x00002_74_q ;
               fgallag0x00003_38 =  fgallag0x00002_76_q ;
               fgallag0x00003_39 =  fgallag0x00002_78_q ;
               fgallag0x00003_40 =  fgallag0x00002_80_q ;
               fgallag0x00003_41 =  fgallag0x00002_82_q ;
               fgallag0x00003_42 =  fgallag0x00002_84_q ;
               fgallag0x00003_43 =  fgallag0x00002_86_q ;
              fgallag0x00003_44 = 
          (!fgallag_sel[2]) ? 
                       fgallag0x00002_88_q: 
                       fgallag0x00002_89_q;
               fgallag0x00003_45 =  0;
