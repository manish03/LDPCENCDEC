// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

`default_nettype none
/*
 *-------------------------------------------------------------
 *
 * user_project_wrapper
 *
 * This wrapper enumerates all of the pins available to the
 * user for the user project.
 *
 * An example user project is provided in this wrapper.  The
 * example should be removed and replaced with the actual
 * user project.
 *
 *-------------------------------------------------------------
 */

module user_project_wrapper #(
    parameter BITS = 32
) (
`ifdef USE_POWER_PINS
    inout vdda1,	// User area 1 3.3V supply
    inout vdda2,	// User area 2 3.3V supply
    inout vssa1,	// User area 1 analog ground
    inout vssa2,	// User area 2 analog ground
    inout vccd1,	// User area 1 1.8V supply
    inout vccd2,	// User area 2 1.8v supply
    inout vssd1,	// User area 1 digital ground
    inout vssd2,	// User area 2 digital ground
`endif

    // Wishbone Slave ports (WB MI A)
    input wb_clk_i,
    input wb_rst_i,
    input wbs_stb_i,
    input wbs_cyc_i,
    input wbs_we_i,
    input [3:0] wbs_sel_i,
    input [31:0] wbs_dat_i,
    input [31:0] wbs_adr_i,
    output wbs_ack_o,
    output [31:0] wbs_dat_o,

    // Logic Analyzer Signals
    input  [127:0] la_data_in,
    output [127:0] la_data_out,
    input  [127:0] la_oenb,

    // IOs
    input  [`MPRJ_IO_PADS-1:0] io_in,
    output [`MPRJ_IO_PADS-1:0] io_out,
    output [`MPRJ_IO_PADS-1:0] io_oeb,

    // Analog (direct connection to GPIO pad---use with caution)
    // Note that analog I/O is not available on the 7 lowest-numbered
    // GPIO pads, and so the analog_io indexing is offset from the
    // GPIO indexing by 7 (also upper 2 GPIOs do not have analog_io).
    inout [`MPRJ_IO_PADS-10:0] analog_io,

    // Independent clock (on independent integer divider)
    input   user_clock2,

    // User maskable interrupt signals
    output [2:0] user_irq
);


wire P_inputnoutput;
wire P_input;
wire [15:0] P_in_out_sel;
wire PO_output;

assign la_data_out = 128'b0;

assign P_in_out_sel[0]  = io_in[5+0]  ;
assign P_in_out_sel[1]  = io_in[5+1]  ;
assign P_in_out_sel[2]  = io_in[5+2]  ;
assign P_in_out_sel[3]  = io_in[5+3]  ;
assign P_in_out_sel[4]  = io_in[5+4]  ;
assign P_in_out_sel[5]  = io_in[5+5]  ;
assign P_in_out_sel[6]  = io_in[5+6]  ;
assign P_in_out_sel[7]  = io_in[5+7]  ;
assign P_in_out_sel[8]  = io_in[5+8]  ;
assign P_in_out_sel[9]  = io_in[5+9]  ;
assign P_in_out_sel[10] = io_in[5+10] ;
assign P_in_out_sel[11] = io_in[5+11] ;
assign P_in_out_sel[12] = io_in[5+12] ;
assign P_in_out_sel[13] = io_in[5+13] ;
assign P_in_out_sel[14] = io_in[5+14] ;
assign P_in_out_sel[15] = io_in[5+15] ;

assign P_inputnoutput   = io_in[5+16] ;
assign P_input          = io_in[5+17] ;


assign io_oeb[4:  0]                  = {(5){1'b1}};                       //input pins
assign io_oeb[5+17:  5]               = {(5+17-5+1){1'b1}};                //input pins
assign io_oeb[5+18]                   = 1'b0;                              //output pins
assign io_oeb[`MPRJ_IO_PADS-1:5+18+1] = {(`MPRJ_IO_PADS-(5+18+1)){1'b1}};  //input pins


assign io_out[4:  0]                  = {(5){1'b0}};                       //input pins
assign io_out[5+17:  5]               = {(5+17-5+1){1'b0}};                //input pins;
assign io_out[5+18]                   = PO_output;                         //output pins //23
assign io_out[`MPRJ_IO_PADS-1:5+18+1] = {(`MPRJ_IO_PADS-(5+18+1)){1'b0}};  //input pins



assign analog_io = {(`MPRJ_IO_PADS-9){1'b0}};
assign user_irq = 3'b0;
/*--------------------------------------*/
/* User project is instantiated  here   */
/*--------------------------------------*/

ldpcEncDec mprj (
`ifdef USE_POWER_PINS
	.vccd1(vccd1),	// User area 1 1.8V power
	.vssd1(vssd1),	// User area 1 digital ground
	.vccd2(vccd2),	// User area 1 1.8V power
	.vssd2(vssd2),	// User area 1 digital ground
`endif

    .wb_clk_i(wb_clk_i),
    .wb_rst_i(wb_rst_i),

    // MGMT SoC Wishbone Slave

    .wbs_cyc_i(wbs_cyc_i),
    .wbs_stb_i(wbs_stb_i),
    .wbs_we_i(wbs_we_i),
    .wbs_sel_i(wbs_sel_i),
    .wbs_adr_i(wbs_adr_i),
    .wbs_dat_i(wbs_dat_i),
    .wbs_ack_o(wbs_ack_o),
    .wbs_dat_o(wbs_dat_o),

    .P_inputnoutput(P_inputnoutput),
    .P_input(P_input),
    .P_in_out_sel(P_in_out_sel),
    .PO_output(PO_output)


);

endmodule	// user_project_wrapper

`default_nettype wire
