assign y_nr_in_port[   0] =  o_LDPC_ENC_MSG_IN_0_msg_in;
assign y_nr_in_port[   1] =  o_LDPC_ENC_MSG_IN_1_msg_in;
assign y_nr_in_port[   2] =  o_LDPC_ENC_MSG_IN_2_msg_in;
assign y_nr_in_port[   3] =  o_LDPC_ENC_MSG_IN_3_msg_in;
assign y_nr_in_port[   4] =  o_LDPC_ENC_MSG_IN_4_msg_in;
assign y_nr_in_port[   5] =  o_LDPC_ENC_MSG_IN_5_msg_in;
assign y_nr_in_port[   6] =  o_LDPC_ENC_MSG_IN_6_msg_in;
assign y_nr_in_port[   7] =  o_LDPC_ENC_MSG_IN_7_msg_in;
assign y_nr_in_port[   8] =  o_LDPC_ENC_MSG_IN_8_msg_in;
assign y_nr_in_port[   9] =  o_LDPC_ENC_MSG_IN_9_msg_in;
assign y_nr_in_port[   10] =  o_LDPC_ENC_MSG_IN_10_msg_in;
assign y_nr_in_port[   11] =  o_LDPC_ENC_MSG_IN_11_msg_in;
assign y_nr_in_port[   12] =  o_LDPC_ENC_MSG_IN_12_msg_in;
assign y_nr_in_port[   13] =  o_LDPC_ENC_MSG_IN_13_msg_in;
assign y_nr_in_port[   14] =  o_LDPC_ENC_MSG_IN_14_msg_in;
assign y_nr_in_port[   15] =  o_LDPC_ENC_MSG_IN_15_msg_in;
assign y_nr_in_port[   16] =  o_LDPC_ENC_MSG_IN_16_msg_in;
assign y_nr_in_port[   17] =  o_LDPC_ENC_MSG_IN_17_msg_in;
assign y_nr_in_port[   18] =  o_LDPC_ENC_MSG_IN_18_msg_in;
assign y_nr_in_port[   19] =  o_LDPC_ENC_MSG_IN_19_msg_in;
assign y_nr_in_port[   20] =  o_LDPC_ENC_MSG_IN_20_msg_in;
assign y_nr_in_port[   21] =  o_LDPC_ENC_MSG_IN_21_msg_in;
assign y_nr_in_port[   22] =  o_LDPC_ENC_MSG_IN_22_msg_in;
assign y_nr_in_port[   23] =  o_LDPC_ENC_MSG_IN_23_msg_in;
assign y_nr_in_port[   24] =  o_LDPC_ENC_MSG_IN_24_msg_in;
assign y_nr_in_port[   25] =  o_LDPC_ENC_MSG_IN_25_msg_in;
assign y_nr_in_port[   26] =  o_LDPC_ENC_MSG_IN_26_msg_in;
assign y_nr_in_port[   27] =  o_LDPC_ENC_MSG_IN_27_msg_in;
assign y_nr_in_port[   28] =  o_LDPC_ENC_MSG_IN_28_msg_in;
assign y_nr_in_port[   29] =  o_LDPC_ENC_MSG_IN_29_msg_in;
assign y_nr_in_port[   30] =  o_LDPC_ENC_MSG_IN_30_msg_in;
assign y_nr_in_port[   31] =  o_LDPC_ENC_MSG_IN_31_msg_in;
assign y_nr_in_port[   32] =  o_LDPC_ENC_MSG_IN_32_msg_in;
assign y_nr_in_port[   33] =  o_LDPC_ENC_MSG_IN_33_msg_in;
assign y_nr_in_port[   34] =  o_LDPC_ENC_MSG_IN_34_msg_in;
assign y_nr_in_port[   35] =  o_LDPC_ENC_MSG_IN_35_msg_in;
assign y_nr_in_port[   36] =  o_LDPC_ENC_MSG_IN_36_msg_in;
assign y_nr_in_port[   37] =  o_LDPC_ENC_MSG_IN_37_msg_in;
assign y_nr_in_port[   38] =  o_LDPC_ENC_MSG_IN_38_msg_in;
assign y_nr_in_port[   39] =  o_LDPC_ENC_MSG_IN_39_msg_in;
assign i_LDPC_ENC_CODEWRD_OUT_0_enc_codeword = y_nr_enc[   0] ;
assign i_LDPC_ENC_CODEWRD_OUT_1_enc_codeword = y_nr_enc[   1] ;
assign i_LDPC_ENC_CODEWRD_OUT_2_enc_codeword = y_nr_enc[   2] ;
assign i_LDPC_ENC_CODEWRD_OUT_3_enc_codeword = y_nr_enc[   3] ;
assign i_LDPC_ENC_CODEWRD_OUT_4_enc_codeword = y_nr_enc[   4] ;
assign i_LDPC_ENC_CODEWRD_OUT_5_enc_codeword = y_nr_enc[   5] ;
assign i_LDPC_ENC_CODEWRD_OUT_6_enc_codeword = y_nr_enc[   6] ;
assign i_LDPC_ENC_CODEWRD_OUT_7_enc_codeword = y_nr_enc[   7] ;
assign i_LDPC_ENC_CODEWRD_OUT_8_enc_codeword = y_nr_enc[   8] ;
assign i_LDPC_ENC_CODEWRD_OUT_9_enc_codeword = y_nr_enc[   9] ;
assign i_LDPC_ENC_CODEWRD_OUT_10_enc_codeword = y_nr_enc[   10] ;
assign i_LDPC_ENC_CODEWRD_OUT_11_enc_codeword = y_nr_enc[   11] ;
assign i_LDPC_ENC_CODEWRD_OUT_12_enc_codeword = y_nr_enc[   12] ;
assign i_LDPC_ENC_CODEWRD_OUT_13_enc_codeword = y_nr_enc[   13] ;
assign i_LDPC_ENC_CODEWRD_OUT_14_enc_codeword = y_nr_enc[   14] ;
assign i_LDPC_ENC_CODEWRD_OUT_15_enc_codeword = y_nr_enc[   15] ;
assign i_LDPC_ENC_CODEWRD_OUT_16_enc_codeword = y_nr_enc[   16] ;
assign i_LDPC_ENC_CODEWRD_OUT_17_enc_codeword = y_nr_enc[   17] ;
assign i_LDPC_ENC_CODEWRD_OUT_18_enc_codeword = y_nr_enc[   18] ;
assign i_LDPC_ENC_CODEWRD_OUT_19_enc_codeword = y_nr_enc[   19] ;
assign i_LDPC_ENC_CODEWRD_OUT_20_enc_codeword = y_nr_enc[   20] ;
assign i_LDPC_ENC_CODEWRD_OUT_21_enc_codeword = y_nr_enc[   21] ;
assign i_LDPC_ENC_CODEWRD_OUT_22_enc_codeword = y_nr_enc[   22] ;
assign i_LDPC_ENC_CODEWRD_OUT_23_enc_codeword = y_nr_enc[   23] ;
assign i_LDPC_ENC_CODEWRD_OUT_24_enc_codeword = y_nr_enc[   24] ;
assign i_LDPC_ENC_CODEWRD_OUT_25_enc_codeword = y_nr_enc[   25] ;
assign i_LDPC_ENC_CODEWRD_OUT_26_enc_codeword = y_nr_enc[   26] ;
assign i_LDPC_ENC_CODEWRD_OUT_27_enc_codeword = y_nr_enc[   27] ;
assign i_LDPC_ENC_CODEWRD_OUT_28_enc_codeword = y_nr_enc[   28] ;
assign i_LDPC_ENC_CODEWRD_OUT_29_enc_codeword = y_nr_enc[   29] ;
assign i_LDPC_ENC_CODEWRD_OUT_30_enc_codeword = y_nr_enc[   30] ;
assign i_LDPC_ENC_CODEWRD_OUT_31_enc_codeword = y_nr_enc[   31] ;
assign i_LDPC_ENC_CODEWRD_OUT_32_enc_codeword = y_nr_enc[   32] ;
assign i_LDPC_ENC_CODEWRD_OUT_33_enc_codeword = y_nr_enc[   33] ;
assign i_LDPC_ENC_CODEWRD_OUT_34_enc_codeword = y_nr_enc[   34] ;
assign i_LDPC_ENC_CODEWRD_OUT_35_enc_codeword = y_nr_enc[   35] ;
assign i_LDPC_ENC_CODEWRD_OUT_36_enc_codeword = y_nr_enc[   36] ;
assign i_LDPC_ENC_CODEWRD_OUT_37_enc_codeword = y_nr_enc[   37] ;
assign i_LDPC_ENC_CODEWRD_OUT_38_enc_codeword = y_nr_enc[   38] ;
assign i_LDPC_ENC_CODEWRD_OUT_39_enc_codeword = y_nr_enc[   39] ;
assign i_LDPC_ENC_CODEWRD_OUT_40_enc_codeword = y_nr_enc[   40] ;
assign i_LDPC_ENC_CODEWRD_OUT_41_enc_codeword = y_nr_enc[   41] ;
assign i_LDPC_ENC_CODEWRD_OUT_42_enc_codeword = y_nr_enc[   42] ;
assign i_LDPC_ENC_CODEWRD_OUT_43_enc_codeword = y_nr_enc[   43] ;
assign i_LDPC_ENC_CODEWRD_OUT_44_enc_codeword = y_nr_enc[   44] ;
assign i_LDPC_ENC_CODEWRD_OUT_45_enc_codeword = y_nr_enc[   45] ;
assign i_LDPC_ENC_CODEWRD_OUT_46_enc_codeword = y_nr_enc[   46] ;
assign i_LDPC_ENC_CODEWRD_OUT_47_enc_codeword = y_nr_enc[   47] ;
assign i_LDPC_ENC_CODEWRD_OUT_48_enc_codeword = y_nr_enc[   48] ;
assign i_LDPC_ENC_CODEWRD_OUT_49_enc_codeword = y_nr_enc[   49] ;
assign i_LDPC_ENC_CODEWRD_OUT_50_enc_codeword = y_nr_enc[   50] ;
assign i_LDPC_ENC_CODEWRD_OUT_51_enc_codeword = y_nr_enc[   51] ;
assign i_LDPC_ENC_CODEWRD_OUT_52_enc_codeword = y_nr_enc[   52] ;
assign i_LDPC_ENC_CODEWRD_OUT_53_enc_codeword = y_nr_enc[   53] ;
assign i_LDPC_ENC_CODEWRD_OUT_54_enc_codeword = y_nr_enc[   54] ;
assign i_LDPC_ENC_CODEWRD_OUT_55_enc_codeword = y_nr_enc[   55] ;
assign i_LDPC_ENC_CODEWRD_OUT_56_enc_codeword = y_nr_enc[   56] ;
assign i_LDPC_ENC_CODEWRD_OUT_57_enc_codeword = y_nr_enc[   57] ;
assign i_LDPC_ENC_CODEWRD_OUT_58_enc_codeword = y_nr_enc[   58] ;
assign i_LDPC_ENC_CODEWRD_OUT_59_enc_codeword = y_nr_enc[   59] ;
assign i_LDPC_ENC_CODEWRD_OUT_60_enc_codeword = y_nr_enc[   60] ;
assign i_LDPC_ENC_CODEWRD_OUT_61_enc_codeword = y_nr_enc[   61] ;
assign i_LDPC_ENC_CODEWRD_OUT_62_enc_codeword = y_nr_enc[   62] ;
assign i_LDPC_ENC_CODEWRD_OUT_63_enc_codeword = y_nr_enc[   63] ;
assign i_LDPC_ENC_CODEWRD_OUT_64_enc_codeword = y_nr_enc[   64] ;
assign i_LDPC_ENC_CODEWRD_OUT_65_enc_codeword = y_nr_enc[   65] ;
assign i_LDPC_ENC_CODEWRD_OUT_66_enc_codeword = y_nr_enc[   66] ;
assign i_LDPC_ENC_CODEWRD_OUT_67_enc_codeword = y_nr_enc[   67] ;
assign i_LDPC_ENC_CODEWRD_OUT_68_enc_codeword = y_nr_enc[   68] ;
assign i_LDPC_ENC_CODEWRD_OUT_69_enc_codeword = y_nr_enc[   69] ;
assign i_LDPC_ENC_CODEWRD_OUT_70_enc_codeword = y_nr_enc[   70] ;
assign i_LDPC_ENC_CODEWRD_OUT_71_enc_codeword = y_nr_enc[   71] ;
assign i_LDPC_ENC_CODEWRD_OUT_72_enc_codeword = y_nr_enc[   72] ;
assign i_LDPC_ENC_CODEWRD_OUT_73_enc_codeword = y_nr_enc[   73] ;
assign i_LDPC_ENC_CODEWRD_OUT_74_enc_codeword = y_nr_enc[   74] ;
assign i_LDPC_ENC_CODEWRD_OUT_75_enc_codeword = y_nr_enc[   75] ;
assign i_LDPC_ENC_CODEWRD_OUT_76_enc_codeword = y_nr_enc[   76] ;
assign i_LDPC_ENC_CODEWRD_OUT_77_enc_codeword = y_nr_enc[   77] ;
assign i_LDPC_ENC_CODEWRD_OUT_78_enc_codeword = y_nr_enc[   78] ;
assign i_LDPC_ENC_CODEWRD_OUT_79_enc_codeword = y_nr_enc[   79] ;
assign i_LDPC_ENC_CODEWRD_OUT_80_enc_codeword = y_nr_enc[   80] ;
assign i_LDPC_ENC_CODEWRD_OUT_81_enc_codeword = y_nr_enc[   81] ;
assign i_LDPC_ENC_CODEWRD_OUT_82_enc_codeword = y_nr_enc[   82] ;
assign i_LDPC_ENC_CODEWRD_OUT_83_enc_codeword = y_nr_enc[   83] ;
assign i_LDPC_ENC_CODEWRD_OUT_84_enc_codeword = y_nr_enc[   84] ;
assign i_LDPC_ENC_CODEWRD_OUT_85_enc_codeword = y_nr_enc[   85] ;
assign i_LDPC_ENC_CODEWRD_OUT_86_enc_codeword = y_nr_enc[   86] ;
assign i_LDPC_ENC_CODEWRD_OUT_87_enc_codeword = y_nr_enc[   87] ;
assign i_LDPC_ENC_CODEWRD_OUT_88_enc_codeword = y_nr_enc[   88] ;
assign i_LDPC_ENC_CODEWRD_OUT_89_enc_codeword = y_nr_enc[   89] ;
assign i_LDPC_ENC_CODEWRD_OUT_90_enc_codeword = y_nr_enc[   90] ;
assign i_LDPC_ENC_CODEWRD_OUT_91_enc_codeword = y_nr_enc[   91] ;
assign i_LDPC_ENC_CODEWRD_OUT_92_enc_codeword = y_nr_enc[   92] ;
assign i_LDPC_ENC_CODEWRD_OUT_93_enc_codeword = y_nr_enc[   93] ;
assign i_LDPC_ENC_CODEWRD_OUT_94_enc_codeword = y_nr_enc[   94] ;
assign i_LDPC_ENC_CODEWRD_OUT_95_enc_codeword = y_nr_enc[   95] ;
assign i_LDPC_ENC_CODEWRD_OUT_96_enc_codeword = y_nr_enc[   96] ;
assign i_LDPC_ENC_CODEWRD_OUT_97_enc_codeword = y_nr_enc[   97] ;
assign i_LDPC_ENC_CODEWRD_OUT_98_enc_codeword = y_nr_enc[   98] ;
assign i_LDPC_ENC_CODEWRD_OUT_99_enc_codeword = y_nr_enc[   99] ;
assign i_LDPC_ENC_CODEWRD_OUT_100_enc_codeword = y_nr_enc[   100] ;
assign i_LDPC_ENC_CODEWRD_OUT_101_enc_codeword = y_nr_enc[   101] ;
assign i_LDPC_ENC_CODEWRD_OUT_102_enc_codeword = y_nr_enc[   102] ;
assign i_LDPC_ENC_CODEWRD_OUT_103_enc_codeword = y_nr_enc[   103] ;
assign i_LDPC_ENC_CODEWRD_OUT_104_enc_codeword = y_nr_enc[   104] ;
assign i_LDPC_ENC_CODEWRD_OUT_105_enc_codeword = y_nr_enc[   105] ;
assign i_LDPC_ENC_CODEWRD_OUT_106_enc_codeword = y_nr_enc[   106] ;
assign i_LDPC_ENC_CODEWRD_OUT_107_enc_codeword = y_nr_enc[   107] ;
assign i_LDPC_ENC_CODEWRD_OUT_108_enc_codeword = y_nr_enc[   108] ;
assign i_LDPC_ENC_CODEWRD_OUT_109_enc_codeword = y_nr_enc[   109] ;
assign i_LDPC_ENC_CODEWRD_OUT_110_enc_codeword = y_nr_enc[   110] ;
assign i_LDPC_ENC_CODEWRD_OUT_111_enc_codeword = y_nr_enc[   111] ;
assign i_LDPC_ENC_CODEWRD_OUT_112_enc_codeword = y_nr_enc[   112] ;
assign i_LDPC_ENC_CODEWRD_OUT_113_enc_codeword = y_nr_enc[   113] ;
assign i_LDPC_ENC_CODEWRD_OUT_114_enc_codeword = y_nr_enc[   114] ;
assign i_LDPC_ENC_CODEWRD_OUT_115_enc_codeword = y_nr_enc[   115] ;
assign i_LDPC_ENC_CODEWRD_OUT_116_enc_codeword = y_nr_enc[   116] ;
assign i_LDPC_ENC_CODEWRD_OUT_117_enc_codeword = y_nr_enc[   117] ;
assign i_LDPC_ENC_CODEWRD_OUT_118_enc_codeword = y_nr_enc[   118] ;
assign i_LDPC_ENC_CODEWRD_OUT_119_enc_codeword = y_nr_enc[   119] ;
assign i_LDPC_ENC_CODEWRD_OUT_120_enc_codeword = y_nr_enc[   120] ;
assign i_LDPC_ENC_CODEWRD_OUT_121_enc_codeword = y_nr_enc[   121] ;
assign i_LDPC_ENC_CODEWRD_OUT_122_enc_codeword = y_nr_enc[   122] ;
assign i_LDPC_ENC_CODEWRD_OUT_123_enc_codeword = y_nr_enc[   123] ;
assign i_LDPC_ENC_CODEWRD_OUT_124_enc_codeword = y_nr_enc[   124] ;
assign i_LDPC_ENC_CODEWRD_OUT_125_enc_codeword = y_nr_enc[   125] ;
assign i_LDPC_ENC_CODEWRD_OUT_126_enc_codeword = y_nr_enc[   126] ;
assign i_LDPC_ENC_CODEWRD_OUT_127_enc_codeword = y_nr_enc[   127] ;
assign i_LDPC_ENC_CODEWRD_OUT_128_enc_codeword = y_nr_enc[   128] ;
assign i_LDPC_ENC_CODEWRD_OUT_129_enc_codeword = y_nr_enc[   129] ;
assign i_LDPC_ENC_CODEWRD_OUT_130_enc_codeword = y_nr_enc[   130] ;
assign i_LDPC_ENC_CODEWRD_OUT_131_enc_codeword = y_nr_enc[   131] ;
assign i_LDPC_ENC_CODEWRD_OUT_132_enc_codeword = y_nr_enc[   132] ;
assign i_LDPC_ENC_CODEWRD_OUT_133_enc_codeword = y_nr_enc[   133] ;
assign i_LDPC_ENC_CODEWRD_OUT_134_enc_codeword = y_nr_enc[   134] ;
assign i_LDPC_ENC_CODEWRD_OUT_135_enc_codeword = y_nr_enc[   135] ;
assign i_LDPC_ENC_CODEWRD_OUT_136_enc_codeword = y_nr_enc[   136] ;
assign i_LDPC_ENC_CODEWRD_OUT_137_enc_codeword = y_nr_enc[   137] ;
assign i_LDPC_ENC_CODEWRD_OUT_138_enc_codeword = y_nr_enc[   138] ;
assign i_LDPC_ENC_CODEWRD_OUT_139_enc_codeword = y_nr_enc[   139] ;
assign i_LDPC_ENC_CODEWRD_OUT_140_enc_codeword = y_nr_enc[   140] ;
assign i_LDPC_ENC_CODEWRD_OUT_141_enc_codeword = y_nr_enc[   141] ;
assign i_LDPC_ENC_CODEWRD_OUT_142_enc_codeword = y_nr_enc[   142] ;
assign i_LDPC_ENC_CODEWRD_OUT_143_enc_codeword = y_nr_enc[   143] ;
assign i_LDPC_ENC_CODEWRD_OUT_144_enc_codeword = y_nr_enc[   144] ;
assign i_LDPC_ENC_CODEWRD_OUT_145_enc_codeword = y_nr_enc[   145] ;
assign i_LDPC_ENC_CODEWRD_OUT_146_enc_codeword = y_nr_enc[   146] ;
assign i_LDPC_ENC_CODEWRD_OUT_147_enc_codeword = y_nr_enc[   147] ;
assign i_LDPC_ENC_CODEWRD_OUT_148_enc_codeword = y_nr_enc[   148] ;
assign i_LDPC_ENC_CODEWRD_OUT_149_enc_codeword = y_nr_enc[   149] ;
assign i_LDPC_ENC_CODEWRD_OUT_150_enc_codeword = y_nr_enc[   150] ;
assign i_LDPC_ENC_CODEWRD_OUT_151_enc_codeword = y_nr_enc[   151] ;
assign i_LDPC_ENC_CODEWRD_OUT_152_enc_codeword = y_nr_enc[   152] ;
assign i_LDPC_ENC_CODEWRD_OUT_153_enc_codeword = y_nr_enc[   153] ;
assign i_LDPC_ENC_CODEWRD_OUT_154_enc_codeword = y_nr_enc[   154] ;
assign i_LDPC_ENC_CODEWRD_OUT_155_enc_codeword = y_nr_enc[   155] ;
assign i_LDPC_ENC_CODEWRD_OUT_156_enc_codeword = y_nr_enc[   156] ;
assign i_LDPC_ENC_CODEWRD_OUT_157_enc_codeword = y_nr_enc[   157] ;
assign i_LDPC_ENC_CODEWRD_OUT_158_enc_codeword = y_nr_enc[   158] ;
assign i_LDPC_ENC_CODEWRD_OUT_159_enc_codeword = y_nr_enc[   159] ;
assign i_LDPC_ENC_CODEWRD_OUT_160_enc_codeword = y_nr_enc[   160] ;
assign i_LDPC_ENC_CODEWRD_OUT_161_enc_codeword = y_nr_enc[   161] ;
assign i_LDPC_ENC_CODEWRD_OUT_162_enc_codeword = y_nr_enc[   162] ;
assign i_LDPC_ENC_CODEWRD_OUT_163_enc_codeword = y_nr_enc[   163] ;
assign i_LDPC_ENC_CODEWRD_OUT_164_enc_codeword = y_nr_enc[   164] ;
assign i_LDPC_ENC_CODEWRD_OUT_165_enc_codeword = y_nr_enc[   165] ;
assign i_LDPC_ENC_CODEWRD_OUT_166_enc_codeword = y_nr_enc[   166] ;
assign i_LDPC_ENC_CODEWRD_OUT_167_enc_codeword = y_nr_enc[   167] ;
assign i_LDPC_ENC_CODEWRD_OUT_168_enc_codeword = y_nr_enc[   168] ;
assign i_LDPC_ENC_CODEWRD_OUT_169_enc_codeword = y_nr_enc[   169] ;
assign i_LDPC_ENC_CODEWRD_OUT_170_enc_codeword = y_nr_enc[   170] ;
assign i_LDPC_ENC_CODEWRD_OUT_171_enc_codeword = y_nr_enc[   171] ;
assign i_LDPC_ENC_CODEWRD_OUT_172_enc_codeword = y_nr_enc[   172] ;
assign i_LDPC_ENC_CODEWRD_OUT_173_enc_codeword = y_nr_enc[   173] ;
assign i_LDPC_ENC_CODEWRD_OUT_174_enc_codeword = y_nr_enc[   174] ;
assign i_LDPC_ENC_CODEWRD_OUT_175_enc_codeword = y_nr_enc[   175] ;
assign i_LDPC_ENC_CODEWRD_OUT_176_enc_codeword = y_nr_enc[   176] ;
assign i_LDPC_ENC_CODEWRD_OUT_177_enc_codeword = y_nr_enc[   177] ;
assign i_LDPC_ENC_CODEWRD_OUT_178_enc_codeword = y_nr_enc[   178] ;
assign i_LDPC_ENC_CODEWRD_OUT_179_enc_codeword = y_nr_enc[   179] ;
assign i_LDPC_ENC_CODEWRD_OUT_180_enc_codeword = y_nr_enc[   180] ;
assign i_LDPC_ENC_CODEWRD_OUT_181_enc_codeword = y_nr_enc[   181] ;
assign i_LDPC_ENC_CODEWRD_OUT_182_enc_codeword = y_nr_enc[   182] ;
assign i_LDPC_ENC_CODEWRD_OUT_183_enc_codeword = y_nr_enc[   183] ;
assign i_LDPC_ENC_CODEWRD_OUT_184_enc_codeword = y_nr_enc[   184] ;
assign i_LDPC_ENC_CODEWRD_OUT_185_enc_codeword = y_nr_enc[   185] ;
assign i_LDPC_ENC_CODEWRD_OUT_186_enc_codeword = y_nr_enc[   186] ;
assign i_LDPC_ENC_CODEWRD_OUT_187_enc_codeword = y_nr_enc[   187] ;
assign i_LDPC_ENC_CODEWRD_OUT_188_enc_codeword = y_nr_enc[   188] ;
assign i_LDPC_ENC_CODEWRD_OUT_189_enc_codeword = y_nr_enc[   189] ;
assign i_LDPC_ENC_CODEWRD_OUT_190_enc_codeword = y_nr_enc[   190] ;
assign i_LDPC_ENC_CODEWRD_OUT_191_enc_codeword = y_nr_enc[   191] ;
assign i_LDPC_ENC_CODEWRD_OUT_192_enc_codeword = y_nr_enc[   192] ;
assign i_LDPC_ENC_CODEWRD_OUT_193_enc_codeword = y_nr_enc[   193] ;
assign i_LDPC_ENC_CODEWRD_OUT_194_enc_codeword = y_nr_enc[   194] ;
assign i_LDPC_ENC_CODEWRD_OUT_195_enc_codeword = y_nr_enc[   195] ;
assign i_LDPC_ENC_CODEWRD_OUT_196_enc_codeword = y_nr_enc[   196] ;
assign i_LDPC_ENC_CODEWRD_OUT_197_enc_codeword = y_nr_enc[   197] ;
assign i_LDPC_ENC_CODEWRD_OUT_198_enc_codeword = y_nr_enc[   198] ;
assign i_LDPC_ENC_CODEWRD_OUT_199_enc_codeword = y_nr_enc[   199] ;
assign i_LDPC_ENC_CODEWRD_OUT_200_enc_codeword = y_nr_enc[   200] ;
assign i_LDPC_ENC_CODEWRD_OUT_201_enc_codeword = y_nr_enc[   201] ;
assign i_LDPC_ENC_CODEWRD_OUT_202_enc_codeword = y_nr_enc[   202] ;
assign i_LDPC_ENC_CODEWRD_OUT_203_enc_codeword = y_nr_enc[   203] ;
assign i_LDPC_ENC_CODEWRD_OUT_204_enc_codeword = y_nr_enc[   204] ;
assign i_LDPC_ENC_CODEWRD_OUT_205_enc_codeword = y_nr_enc[   205] ;
assign i_LDPC_ENC_CODEWRD_OUT_206_enc_codeword = y_nr_enc[   206] ;
assign i_LDPC_ENC_CODEWRD_OUT_207_enc_codeword = y_nr_enc[   207] ;
assign i_LDPC_ENC_CODEWRD_VLD_enc_codeword_valid =  valid_cword_enc;
assign sel_q0_0_frmC =  o_LDPC_DEC_SEL_Q0_0_FRMC_sel_q0_0_frmC;
assign sel_q0_1_frmC =  o_LDPC_DEC_SEL_Q0_1_FRMC_sel_q0_1_frmC;
assign err_intro_q0_0_frmC[0] =  o_LDPC_DEC_ERR_Q0_0_INTRO_0_err_intro_q0_0_0;
assign err_intro_q0_0_frmC[1] =  o_LDPC_DEC_ERR_Q0_0_INTRO_1_err_intro_q0_0_1;
assign err_intro_q0_0_frmC[2] =  o_LDPC_DEC_ERR_Q0_0_INTRO_2_err_intro_q0_0_2;
assign err_intro_q0_0_frmC[3] =  o_LDPC_DEC_ERR_Q0_0_INTRO_3_err_intro_q0_0_3;
assign err_intro_q0_0_frmC[4] =  o_LDPC_DEC_ERR_Q0_0_INTRO_4_err_intro_q0_0_4;
assign err_intro_q0_0_frmC[5] =  o_LDPC_DEC_ERR_Q0_0_INTRO_5_err_intro_q0_0_5;
assign err_intro_q0_0_frmC[6] =  o_LDPC_DEC_ERR_Q0_0_INTRO_6_err_intro_q0_0_6;
assign err_intro_q0_0_frmC[7] =  o_LDPC_DEC_ERR_Q0_0_INTRO_7_err_intro_q0_0_7;
assign err_intro_q0_0_frmC[8] =  o_LDPC_DEC_ERR_Q0_0_INTRO_8_err_intro_q0_0_8;
assign err_intro_q0_0_frmC[9] =  o_LDPC_DEC_ERR_Q0_0_INTRO_9_err_intro_q0_0_9;
assign err_intro_q0_0_frmC[10] =  o_LDPC_DEC_ERR_Q0_0_INTRO_10_err_intro_q0_0_10;
assign err_intro_q0_0_frmC[11] =  o_LDPC_DEC_ERR_Q0_0_INTRO_11_err_intro_q0_0_11;
assign err_intro_q0_0_frmC[12] =  o_LDPC_DEC_ERR_Q0_0_INTRO_12_err_intro_q0_0_12;
assign err_intro_q0_0_frmC[13] =  o_LDPC_DEC_ERR_Q0_0_INTRO_13_err_intro_q0_0_13;
assign err_intro_q0_0_frmC[14] =  o_LDPC_DEC_ERR_Q0_0_INTRO_14_err_intro_q0_0_14;
assign err_intro_q0_0_frmC[15] =  o_LDPC_DEC_ERR_Q0_0_INTRO_15_err_intro_q0_0_15;
assign err_intro_q0_0_frmC[16] =  o_LDPC_DEC_ERR_Q0_0_INTRO_16_err_intro_q0_0_16;
assign err_intro_q0_0_frmC[17] =  o_LDPC_DEC_ERR_Q0_0_INTRO_17_err_intro_q0_0_17;
assign err_intro_q0_0_frmC[18] =  o_LDPC_DEC_ERR_Q0_0_INTRO_18_err_intro_q0_0_18;
assign err_intro_q0_0_frmC[19] =  o_LDPC_DEC_ERR_Q0_0_INTRO_19_err_intro_q0_0_19;
assign err_intro_q0_0_frmC[20] =  o_LDPC_DEC_ERR_Q0_0_INTRO_20_err_intro_q0_0_20;
assign err_intro_q0_0_frmC[21] =  o_LDPC_DEC_ERR_Q0_0_INTRO_21_err_intro_q0_0_21;
assign err_intro_q0_0_frmC[22] =  o_LDPC_DEC_ERR_Q0_0_INTRO_22_err_intro_q0_0_22;
assign err_intro_q0_0_frmC[23] =  o_LDPC_DEC_ERR_Q0_0_INTRO_23_err_intro_q0_0_23;
assign err_intro_q0_0_frmC[24] =  o_LDPC_DEC_ERR_Q0_0_INTRO_24_err_intro_q0_0_24;
assign err_intro_q0_0_frmC[25] =  o_LDPC_DEC_ERR_Q0_0_INTRO_25_err_intro_q0_0_25;
assign err_intro_q0_0_frmC[26] =  o_LDPC_DEC_ERR_Q0_0_INTRO_26_err_intro_q0_0_26;
assign err_intro_q0_0_frmC[27] =  o_LDPC_DEC_ERR_Q0_0_INTRO_27_err_intro_q0_0_27;
assign err_intro_q0_0_frmC[28] =  o_LDPC_DEC_ERR_Q0_0_INTRO_28_err_intro_q0_0_28;
assign err_intro_q0_0_frmC[29] =  o_LDPC_DEC_ERR_Q0_0_INTRO_29_err_intro_q0_0_29;
assign err_intro_q0_0_frmC[30] =  o_LDPC_DEC_ERR_Q0_0_INTRO_30_err_intro_q0_0_30;
assign err_intro_q0_0_frmC[31] =  o_LDPC_DEC_ERR_Q0_0_INTRO_31_err_intro_q0_0_31;
assign err_intro_q0_0_frmC[32] =  o_LDPC_DEC_ERR_Q0_0_INTRO_32_err_intro_q0_0_32;
assign err_intro_q0_0_frmC[33] =  o_LDPC_DEC_ERR_Q0_0_INTRO_33_err_intro_q0_0_33;
assign err_intro_q0_0_frmC[34] =  o_LDPC_DEC_ERR_Q0_0_INTRO_34_err_intro_q0_0_34;
assign err_intro_q0_0_frmC[35] =  o_LDPC_DEC_ERR_Q0_0_INTRO_35_err_intro_q0_0_35;
assign err_intro_q0_0_frmC[36] =  o_LDPC_DEC_ERR_Q0_0_INTRO_36_err_intro_q0_0_36;
assign err_intro_q0_0_frmC[37] =  o_LDPC_DEC_ERR_Q0_0_INTRO_37_err_intro_q0_0_37;
assign err_intro_q0_0_frmC[38] =  o_LDPC_DEC_ERR_Q0_0_INTRO_38_err_intro_q0_0_38;
assign err_intro_q0_0_frmC[39] =  o_LDPC_DEC_ERR_Q0_0_INTRO_39_err_intro_q0_0_39;
assign err_intro_q0_0_frmC[40] =  o_LDPC_DEC_ERR_Q0_0_INTRO_40_err_intro_q0_0_40;
assign err_intro_q0_0_frmC[41] =  o_LDPC_DEC_ERR_Q0_0_INTRO_41_err_intro_q0_0_41;
assign err_intro_q0_0_frmC[42] =  o_LDPC_DEC_ERR_Q0_0_INTRO_42_err_intro_q0_0_42;
assign err_intro_q0_0_frmC[43] =  o_LDPC_DEC_ERR_Q0_0_INTRO_43_err_intro_q0_0_43;
assign err_intro_q0_0_frmC[44] =  o_LDPC_DEC_ERR_Q0_0_INTRO_44_err_intro_q0_0_44;
assign err_intro_q0_0_frmC[45] =  o_LDPC_DEC_ERR_Q0_0_INTRO_45_err_intro_q0_0_45;
assign err_intro_q0_0_frmC[46] =  o_LDPC_DEC_ERR_Q0_0_INTRO_46_err_intro_q0_0_46;
assign err_intro_q0_0_frmC[47] =  o_LDPC_DEC_ERR_Q0_0_INTRO_47_err_intro_q0_0_47;
assign err_intro_q0_0_frmC[48] =  o_LDPC_DEC_ERR_Q0_0_INTRO_48_err_intro_q0_0_48;
assign err_intro_q0_0_frmC[49] =  o_LDPC_DEC_ERR_Q0_0_INTRO_49_err_intro_q0_0_49;
assign err_intro_q0_0_frmC[50] =  o_LDPC_DEC_ERR_Q0_0_INTRO_50_err_intro_q0_0_50;
assign err_intro_q0_0_frmC[51] =  o_LDPC_DEC_ERR_Q0_0_INTRO_51_err_intro_q0_0_51;
assign err_intro_q0_0_frmC[52] =  o_LDPC_DEC_ERR_Q0_0_INTRO_52_err_intro_q0_0_52;
assign err_intro_q0_0_frmC[53] =  o_LDPC_DEC_ERR_Q0_0_INTRO_53_err_intro_q0_0_53;
assign err_intro_q0_0_frmC[54] =  o_LDPC_DEC_ERR_Q0_0_INTRO_54_err_intro_q0_0_54;
assign err_intro_q0_0_frmC[55] =  o_LDPC_DEC_ERR_Q0_0_INTRO_55_err_intro_q0_0_55;
assign err_intro_q0_0_frmC[56] =  o_LDPC_DEC_ERR_Q0_0_INTRO_56_err_intro_q0_0_56;
assign err_intro_q0_0_frmC[57] =  o_LDPC_DEC_ERR_Q0_0_INTRO_57_err_intro_q0_0_57;
assign err_intro_q0_0_frmC[58] =  o_LDPC_DEC_ERR_Q0_0_INTRO_58_err_intro_q0_0_58;
assign err_intro_q0_0_frmC[59] =  o_LDPC_DEC_ERR_Q0_0_INTRO_59_err_intro_q0_0_59;
assign err_intro_q0_0_frmC[60] =  o_LDPC_DEC_ERR_Q0_0_INTRO_60_err_intro_q0_0_60;
assign err_intro_q0_0_frmC[61] =  o_LDPC_DEC_ERR_Q0_0_INTRO_61_err_intro_q0_0_61;
assign err_intro_q0_0_frmC[62] =  o_LDPC_DEC_ERR_Q0_0_INTRO_62_err_intro_q0_0_62;
assign err_intro_q0_0_frmC[63] =  o_LDPC_DEC_ERR_Q0_0_INTRO_63_err_intro_q0_0_63;
assign err_intro_q0_0_frmC[64] =  o_LDPC_DEC_ERR_Q0_0_INTRO_64_err_intro_q0_0_64;
assign err_intro_q0_0_frmC[65] =  o_LDPC_DEC_ERR_Q0_0_INTRO_65_err_intro_q0_0_65;
assign err_intro_q0_0_frmC[66] =  o_LDPC_DEC_ERR_Q0_0_INTRO_66_err_intro_q0_0_66;
assign err_intro_q0_0_frmC[67] =  o_LDPC_DEC_ERR_Q0_0_INTRO_67_err_intro_q0_0_67;
assign err_intro_q0_0_frmC[68] =  o_LDPC_DEC_ERR_Q0_0_INTRO_68_err_intro_q0_0_68;
assign err_intro_q0_0_frmC[69] =  o_LDPC_DEC_ERR_Q0_0_INTRO_69_err_intro_q0_0_69;
assign err_intro_q0_0_frmC[70] =  o_LDPC_DEC_ERR_Q0_0_INTRO_70_err_intro_q0_0_70;
assign err_intro_q0_0_frmC[71] =  o_LDPC_DEC_ERR_Q0_0_INTRO_71_err_intro_q0_0_71;
assign err_intro_q0_0_frmC[72] =  o_LDPC_DEC_ERR_Q0_0_INTRO_72_err_intro_q0_0_72;
assign err_intro_q0_0_frmC[73] =  o_LDPC_DEC_ERR_Q0_0_INTRO_73_err_intro_q0_0_73;
assign err_intro_q0_0_frmC[74] =  o_LDPC_DEC_ERR_Q0_0_INTRO_74_err_intro_q0_0_74;
assign err_intro_q0_0_frmC[75] =  o_LDPC_DEC_ERR_Q0_0_INTRO_75_err_intro_q0_0_75;
assign err_intro_q0_0_frmC[76] =  o_LDPC_DEC_ERR_Q0_0_INTRO_76_err_intro_q0_0_76;
assign err_intro_q0_0_frmC[77] =  o_LDPC_DEC_ERR_Q0_0_INTRO_77_err_intro_q0_0_77;
assign err_intro_q0_0_frmC[78] =  o_LDPC_DEC_ERR_Q0_0_INTRO_78_err_intro_q0_0_78;
assign err_intro_q0_0_frmC[79] =  o_LDPC_DEC_ERR_Q0_0_INTRO_79_err_intro_q0_0_79;
assign err_intro_q0_0_frmC[80] =  o_LDPC_DEC_ERR_Q0_0_INTRO_80_err_intro_q0_0_80;
assign err_intro_q0_0_frmC[81] =  o_LDPC_DEC_ERR_Q0_0_INTRO_81_err_intro_q0_0_81;
assign err_intro_q0_0_frmC[82] =  o_LDPC_DEC_ERR_Q0_0_INTRO_82_err_intro_q0_0_82;
assign err_intro_q0_0_frmC[83] =  o_LDPC_DEC_ERR_Q0_0_INTRO_83_err_intro_q0_0_83;
assign err_intro_q0_0_frmC[84] =  o_LDPC_DEC_ERR_Q0_0_INTRO_84_err_intro_q0_0_84;
assign err_intro_q0_0_frmC[85] =  o_LDPC_DEC_ERR_Q0_0_INTRO_85_err_intro_q0_0_85;
assign err_intro_q0_0_frmC[86] =  o_LDPC_DEC_ERR_Q0_0_INTRO_86_err_intro_q0_0_86;
assign err_intro_q0_0_frmC[87] =  o_LDPC_DEC_ERR_Q0_0_INTRO_87_err_intro_q0_0_87;
assign err_intro_q0_0_frmC[88] =  o_LDPC_DEC_ERR_Q0_0_INTRO_88_err_intro_q0_0_88;
assign err_intro_q0_0_frmC[89] =  o_LDPC_DEC_ERR_Q0_0_INTRO_89_err_intro_q0_0_89;
assign err_intro_q0_0_frmC[90] =  o_LDPC_DEC_ERR_Q0_0_INTRO_90_err_intro_q0_0_90;
assign err_intro_q0_0_frmC[91] =  o_LDPC_DEC_ERR_Q0_0_INTRO_91_err_intro_q0_0_91;
assign err_intro_q0_0_frmC[92] =  o_LDPC_DEC_ERR_Q0_0_INTRO_92_err_intro_q0_0_92;
assign err_intro_q0_0_frmC[93] =  o_LDPC_DEC_ERR_Q0_0_INTRO_93_err_intro_q0_0_93;
assign err_intro_q0_0_frmC[94] =  o_LDPC_DEC_ERR_Q0_0_INTRO_94_err_intro_q0_0_94;
assign err_intro_q0_0_frmC[95] =  o_LDPC_DEC_ERR_Q0_0_INTRO_95_err_intro_q0_0_95;
assign err_intro_q0_0_frmC[96] =  o_LDPC_DEC_ERR_Q0_0_INTRO_96_err_intro_q0_0_96;
assign err_intro_q0_0_frmC[97] =  o_LDPC_DEC_ERR_Q0_0_INTRO_97_err_intro_q0_0_97;
assign err_intro_q0_0_frmC[98] =  o_LDPC_DEC_ERR_Q0_0_INTRO_98_err_intro_q0_0_98;
assign err_intro_q0_0_frmC[99] =  o_LDPC_DEC_ERR_Q0_0_INTRO_99_err_intro_q0_0_99;
assign err_intro_q0_0_frmC[100] =  o_LDPC_DEC_ERR_Q0_0_INTRO_100_err_intro_q0_0_100;
assign err_intro_q0_0_frmC[101] =  o_LDPC_DEC_ERR_Q0_0_INTRO_101_err_intro_q0_0_101;
assign err_intro_q0_0_frmC[102] =  o_LDPC_DEC_ERR_Q0_0_INTRO_102_err_intro_q0_0_102;
assign err_intro_q0_0_frmC[103] =  o_LDPC_DEC_ERR_Q0_0_INTRO_103_err_intro_q0_0_103;
assign err_intro_q0_0_frmC[104] =  o_LDPC_DEC_ERR_Q0_0_INTRO_104_err_intro_q0_0_104;
assign err_intro_q0_0_frmC[105] =  o_LDPC_DEC_ERR_Q0_0_INTRO_105_err_intro_q0_0_105;
assign err_intro_q0_0_frmC[106] =  o_LDPC_DEC_ERR_Q0_0_INTRO_106_err_intro_q0_0_106;
assign err_intro_q0_0_frmC[107] =  o_LDPC_DEC_ERR_Q0_0_INTRO_107_err_intro_q0_0_107;
assign err_intro_q0_0_frmC[108] =  o_LDPC_DEC_ERR_Q0_0_INTRO_108_err_intro_q0_0_108;
assign err_intro_q0_0_frmC[109] =  o_LDPC_DEC_ERR_Q0_0_INTRO_109_err_intro_q0_0_109;
assign err_intro_q0_0_frmC[110] =  o_LDPC_DEC_ERR_Q0_0_INTRO_110_err_intro_q0_0_110;
assign err_intro_q0_0_frmC[111] =  o_LDPC_DEC_ERR_Q0_0_INTRO_111_err_intro_q0_0_111;
assign err_intro_q0_0_frmC[112] =  o_LDPC_DEC_ERR_Q0_0_INTRO_112_err_intro_q0_0_112;
assign err_intro_q0_0_frmC[113] =  o_LDPC_DEC_ERR_Q0_0_INTRO_113_err_intro_q0_0_113;
assign err_intro_q0_0_frmC[114] =  o_LDPC_DEC_ERR_Q0_0_INTRO_114_err_intro_q0_0_114;
assign err_intro_q0_0_frmC[115] =  o_LDPC_DEC_ERR_Q0_0_INTRO_115_err_intro_q0_0_115;
assign err_intro_q0_0_frmC[116] =  o_LDPC_DEC_ERR_Q0_0_INTRO_116_err_intro_q0_0_116;
assign err_intro_q0_0_frmC[117] =  o_LDPC_DEC_ERR_Q0_0_INTRO_117_err_intro_q0_0_117;
assign err_intro_q0_0_frmC[118] =  o_LDPC_DEC_ERR_Q0_0_INTRO_118_err_intro_q0_0_118;
assign err_intro_q0_0_frmC[119] =  o_LDPC_DEC_ERR_Q0_0_INTRO_119_err_intro_q0_0_119;
assign err_intro_q0_0_frmC[120] =  o_LDPC_DEC_ERR_Q0_0_INTRO_120_err_intro_q0_0_120;
assign err_intro_q0_0_frmC[121] =  o_LDPC_DEC_ERR_Q0_0_INTRO_121_err_intro_q0_0_121;
assign err_intro_q0_0_frmC[122] =  o_LDPC_DEC_ERR_Q0_0_INTRO_122_err_intro_q0_0_122;
assign err_intro_q0_0_frmC[123] =  o_LDPC_DEC_ERR_Q0_0_INTRO_123_err_intro_q0_0_123;
assign err_intro_q0_0_frmC[124] =  o_LDPC_DEC_ERR_Q0_0_INTRO_124_err_intro_q0_0_124;
assign err_intro_q0_0_frmC[125] =  o_LDPC_DEC_ERR_Q0_0_INTRO_125_err_intro_q0_0_125;
assign err_intro_q0_0_frmC[126] =  o_LDPC_DEC_ERR_Q0_0_INTRO_126_err_intro_q0_0_126;
assign err_intro_q0_0_frmC[127] =  o_LDPC_DEC_ERR_Q0_0_INTRO_127_err_intro_q0_0_127;
assign err_intro_q0_0_frmC[128] =  o_LDPC_DEC_ERR_Q0_0_INTRO_128_err_intro_q0_0_128;
assign err_intro_q0_0_frmC[129] =  o_LDPC_DEC_ERR_Q0_0_INTRO_129_err_intro_q0_0_129;
assign err_intro_q0_0_frmC[130] =  o_LDPC_DEC_ERR_Q0_0_INTRO_130_err_intro_q0_0_130;
assign err_intro_q0_0_frmC[131] =  o_LDPC_DEC_ERR_Q0_0_INTRO_131_err_intro_q0_0_131;
assign err_intro_q0_0_frmC[132] =  o_LDPC_DEC_ERR_Q0_0_INTRO_132_err_intro_q0_0_132;
assign err_intro_q0_0_frmC[133] =  o_LDPC_DEC_ERR_Q0_0_INTRO_133_err_intro_q0_0_133;
assign err_intro_q0_0_frmC[134] =  o_LDPC_DEC_ERR_Q0_0_INTRO_134_err_intro_q0_0_134;
assign err_intro_q0_0_frmC[135] =  o_LDPC_DEC_ERR_Q0_0_INTRO_135_err_intro_q0_0_135;
assign err_intro_q0_0_frmC[136] =  o_LDPC_DEC_ERR_Q0_0_INTRO_136_err_intro_q0_0_136;
assign err_intro_q0_0_frmC[137] =  o_LDPC_DEC_ERR_Q0_0_INTRO_137_err_intro_q0_0_137;
assign err_intro_q0_0_frmC[138] =  o_LDPC_DEC_ERR_Q0_0_INTRO_138_err_intro_q0_0_138;
assign err_intro_q0_0_frmC[139] =  o_LDPC_DEC_ERR_Q0_0_INTRO_139_err_intro_q0_0_139;
assign err_intro_q0_0_frmC[140] =  o_LDPC_DEC_ERR_Q0_0_INTRO_140_err_intro_q0_0_140;
assign err_intro_q0_0_frmC[141] =  o_LDPC_DEC_ERR_Q0_0_INTRO_141_err_intro_q0_0_141;
assign err_intro_q0_0_frmC[142] =  o_LDPC_DEC_ERR_Q0_0_INTRO_142_err_intro_q0_0_142;
assign err_intro_q0_0_frmC[143] =  o_LDPC_DEC_ERR_Q0_0_INTRO_143_err_intro_q0_0_143;
assign err_intro_q0_0_frmC[144] =  o_LDPC_DEC_ERR_Q0_0_INTRO_144_err_intro_q0_0_144;
assign err_intro_q0_0_frmC[145] =  o_LDPC_DEC_ERR_Q0_0_INTRO_145_err_intro_q0_0_145;
assign err_intro_q0_0_frmC[146] =  o_LDPC_DEC_ERR_Q0_0_INTRO_146_err_intro_q0_0_146;
assign err_intro_q0_0_frmC[147] =  o_LDPC_DEC_ERR_Q0_0_INTRO_147_err_intro_q0_0_147;
assign err_intro_q0_0_frmC[148] =  o_LDPC_DEC_ERR_Q0_0_INTRO_148_err_intro_q0_0_148;
assign err_intro_q0_0_frmC[149] =  o_LDPC_DEC_ERR_Q0_0_INTRO_149_err_intro_q0_0_149;
assign err_intro_q0_0_frmC[150] =  o_LDPC_DEC_ERR_Q0_0_INTRO_150_err_intro_q0_0_150;
assign err_intro_q0_0_frmC[151] =  o_LDPC_DEC_ERR_Q0_0_INTRO_151_err_intro_q0_0_151;
assign err_intro_q0_0_frmC[152] =  o_LDPC_DEC_ERR_Q0_0_INTRO_152_err_intro_q0_0_152;
assign err_intro_q0_0_frmC[153] =  o_LDPC_DEC_ERR_Q0_0_INTRO_153_err_intro_q0_0_153;
assign err_intro_q0_0_frmC[154] =  o_LDPC_DEC_ERR_Q0_0_INTRO_154_err_intro_q0_0_154;
assign err_intro_q0_0_frmC[155] =  o_LDPC_DEC_ERR_Q0_0_INTRO_155_err_intro_q0_0_155;
assign err_intro_q0_0_frmC[156] =  o_LDPC_DEC_ERR_Q0_0_INTRO_156_err_intro_q0_0_156;
assign err_intro_q0_0_frmC[157] =  o_LDPC_DEC_ERR_Q0_0_INTRO_157_err_intro_q0_0_157;
assign err_intro_q0_0_frmC[158] =  o_LDPC_DEC_ERR_Q0_0_INTRO_158_err_intro_q0_0_158;
assign err_intro_q0_0_frmC[159] =  o_LDPC_DEC_ERR_Q0_0_INTRO_159_err_intro_q0_0_159;
assign err_intro_q0_0_frmC[160] =  o_LDPC_DEC_ERR_Q0_0_INTRO_160_err_intro_q0_0_160;
assign err_intro_q0_0_frmC[161] =  o_LDPC_DEC_ERR_Q0_0_INTRO_161_err_intro_q0_0_161;
assign err_intro_q0_0_frmC[162] =  o_LDPC_DEC_ERR_Q0_0_INTRO_162_err_intro_q0_0_162;
assign err_intro_q0_0_frmC[163] =  o_LDPC_DEC_ERR_Q0_0_INTRO_163_err_intro_q0_0_163;
assign err_intro_q0_0_frmC[164] =  o_LDPC_DEC_ERR_Q0_0_INTRO_164_err_intro_q0_0_164;
assign err_intro_q0_0_frmC[165] =  o_LDPC_DEC_ERR_Q0_0_INTRO_165_err_intro_q0_0_165;
assign err_intro_q0_0_frmC[166] =  o_LDPC_DEC_ERR_Q0_0_INTRO_166_err_intro_q0_0_166;
assign err_intro_q0_0_frmC[167] =  o_LDPC_DEC_ERR_Q0_0_INTRO_167_err_intro_q0_0_167;
assign err_intro_q0_0_frmC[168] =  o_LDPC_DEC_ERR_Q0_0_INTRO_168_err_intro_q0_0_168;
assign err_intro_q0_0_frmC[169] =  o_LDPC_DEC_ERR_Q0_0_INTRO_169_err_intro_q0_0_169;
assign err_intro_q0_0_frmC[170] =  o_LDPC_DEC_ERR_Q0_0_INTRO_170_err_intro_q0_0_170;
assign err_intro_q0_0_frmC[171] =  o_LDPC_DEC_ERR_Q0_0_INTRO_171_err_intro_q0_0_171;
assign err_intro_q0_0_frmC[172] =  o_LDPC_DEC_ERR_Q0_0_INTRO_172_err_intro_q0_0_172;
assign err_intro_q0_0_frmC[173] =  o_LDPC_DEC_ERR_Q0_0_INTRO_173_err_intro_q0_0_173;
assign err_intro_q0_0_frmC[174] =  o_LDPC_DEC_ERR_Q0_0_INTRO_174_err_intro_q0_0_174;
assign err_intro_q0_0_frmC[175] =  o_LDPC_DEC_ERR_Q0_0_INTRO_175_err_intro_q0_0_175;
assign err_intro_q0_0_frmC[176] =  o_LDPC_DEC_ERR_Q0_0_INTRO_176_err_intro_q0_0_176;
assign err_intro_q0_0_frmC[177] =  o_LDPC_DEC_ERR_Q0_0_INTRO_177_err_intro_q0_0_177;
assign err_intro_q0_0_frmC[178] =  o_LDPC_DEC_ERR_Q0_0_INTRO_178_err_intro_q0_0_178;
assign err_intro_q0_0_frmC[179] =  o_LDPC_DEC_ERR_Q0_0_INTRO_179_err_intro_q0_0_179;
assign err_intro_q0_0_frmC[180] =  o_LDPC_DEC_ERR_Q0_0_INTRO_180_err_intro_q0_0_180;
assign err_intro_q0_0_frmC[181] =  o_LDPC_DEC_ERR_Q0_0_INTRO_181_err_intro_q0_0_181;
assign err_intro_q0_0_frmC[182] =  o_LDPC_DEC_ERR_Q0_0_INTRO_182_err_intro_q0_0_182;
assign err_intro_q0_0_frmC[183] =  o_LDPC_DEC_ERR_Q0_0_INTRO_183_err_intro_q0_0_183;
assign err_intro_q0_0_frmC[184] =  o_LDPC_DEC_ERR_Q0_0_INTRO_184_err_intro_q0_0_184;
assign err_intro_q0_0_frmC[185] =  o_LDPC_DEC_ERR_Q0_0_INTRO_185_err_intro_q0_0_185;
assign err_intro_q0_0_frmC[186] =  o_LDPC_DEC_ERR_Q0_0_INTRO_186_err_intro_q0_0_186;
assign err_intro_q0_0_frmC[187] =  o_LDPC_DEC_ERR_Q0_0_INTRO_187_err_intro_q0_0_187;
assign err_intro_q0_0_frmC[188] =  o_LDPC_DEC_ERR_Q0_0_INTRO_188_err_intro_q0_0_188;
assign err_intro_q0_0_frmC[189] =  o_LDPC_DEC_ERR_Q0_0_INTRO_189_err_intro_q0_0_189;
assign err_intro_q0_0_frmC[190] =  o_LDPC_DEC_ERR_Q0_0_INTRO_190_err_intro_q0_0_190;
assign err_intro_q0_0_frmC[191] =  o_LDPC_DEC_ERR_Q0_0_INTRO_191_err_intro_q0_0_191;
assign err_intro_q0_0_frmC[192] =  o_LDPC_DEC_ERR_Q0_0_INTRO_192_err_intro_q0_0_192;
assign err_intro_q0_0_frmC[193] =  o_LDPC_DEC_ERR_Q0_0_INTRO_193_err_intro_q0_0_193;
assign err_intro_q0_0_frmC[194] =  o_LDPC_DEC_ERR_Q0_0_INTRO_194_err_intro_q0_0_194;
assign err_intro_q0_0_frmC[195] =  o_LDPC_DEC_ERR_Q0_0_INTRO_195_err_intro_q0_0_195;
assign err_intro_q0_0_frmC[196] =  o_LDPC_DEC_ERR_Q0_0_INTRO_196_err_intro_q0_0_196;
assign err_intro_q0_0_frmC[197] =  o_LDPC_DEC_ERR_Q0_0_INTRO_197_err_intro_q0_0_197;
assign err_intro_q0_0_frmC[198] =  o_LDPC_DEC_ERR_Q0_0_INTRO_198_err_intro_q0_0_198;
assign err_intro_q0_0_frmC[199] =  o_LDPC_DEC_ERR_Q0_0_INTRO_199_err_intro_q0_0_199;
assign err_intro_q0_0_frmC[200] =  o_LDPC_DEC_ERR_Q0_0_INTRO_200_err_intro_q0_0_200;
assign err_intro_q0_0_frmC[201] =  o_LDPC_DEC_ERR_Q0_0_INTRO_201_err_intro_q0_0_201;
assign err_intro_q0_0_frmC[202] =  o_LDPC_DEC_ERR_Q0_0_INTRO_202_err_intro_q0_0_202;
assign err_intro_q0_0_frmC[203] =  o_LDPC_DEC_ERR_Q0_0_INTRO_203_err_intro_q0_0_203;
assign err_intro_q0_0_frmC[204] =  o_LDPC_DEC_ERR_Q0_0_INTRO_204_err_intro_q0_0_204;
assign err_intro_q0_0_frmC[205] =  o_LDPC_DEC_ERR_Q0_0_INTRO_205_err_intro_q0_0_205;
assign err_intro_q0_0_frmC[206] =  o_LDPC_DEC_ERR_Q0_0_INTRO_206_err_intro_q0_0_206;
assign err_intro_q0_0_frmC[207] =  o_LDPC_DEC_ERR_Q0_0_INTRO_207_err_intro_q0_0_207;
assign err_intro_q0_1_frmC[0] =  o_LDPC_DEC_ERR_Q0_1_INTRO_0_err_intro_q0_1_0;
assign err_intro_q0_1_frmC[1] =  o_LDPC_DEC_ERR_Q0_1_INTRO_1_err_intro_q0_1_1;
assign err_intro_q0_1_frmC[2] =  o_LDPC_DEC_ERR_Q0_1_INTRO_2_err_intro_q0_1_2;
assign err_intro_q0_1_frmC[3] =  o_LDPC_DEC_ERR_Q0_1_INTRO_3_err_intro_q0_1_3;
assign err_intro_q0_1_frmC[4] =  o_LDPC_DEC_ERR_Q0_1_INTRO_4_err_intro_q0_1_4;
assign err_intro_q0_1_frmC[5] =  o_LDPC_DEC_ERR_Q0_1_INTRO_5_err_intro_q0_1_5;
assign err_intro_q0_1_frmC[6] =  o_LDPC_DEC_ERR_Q0_1_INTRO_6_err_intro_q0_1_6;
assign err_intro_q0_1_frmC[7] =  o_LDPC_DEC_ERR_Q0_1_INTRO_7_err_intro_q0_1_7;
assign err_intro_q0_1_frmC[8] =  o_LDPC_DEC_ERR_Q0_1_INTRO_8_err_intro_q0_1_8;
assign err_intro_q0_1_frmC[9] =  o_LDPC_DEC_ERR_Q0_1_INTRO_9_err_intro_q0_1_9;
assign err_intro_q0_1_frmC[10] =  o_LDPC_DEC_ERR_Q0_1_INTRO_10_err_intro_q0_1_10;
assign err_intro_q0_1_frmC[11] =  o_LDPC_DEC_ERR_Q0_1_INTRO_11_err_intro_q0_1_11;
assign err_intro_q0_1_frmC[12] =  o_LDPC_DEC_ERR_Q0_1_INTRO_12_err_intro_q0_1_12;
assign err_intro_q0_1_frmC[13] =  o_LDPC_DEC_ERR_Q0_1_INTRO_13_err_intro_q0_1_13;
assign err_intro_q0_1_frmC[14] =  o_LDPC_DEC_ERR_Q0_1_INTRO_14_err_intro_q0_1_14;
assign err_intro_q0_1_frmC[15] =  o_LDPC_DEC_ERR_Q0_1_INTRO_15_err_intro_q0_1_15;
assign err_intro_q0_1_frmC[16] =  o_LDPC_DEC_ERR_Q0_1_INTRO_16_err_intro_q0_1_16;
assign err_intro_q0_1_frmC[17] =  o_LDPC_DEC_ERR_Q0_1_INTRO_17_err_intro_q0_1_17;
assign err_intro_q0_1_frmC[18] =  o_LDPC_DEC_ERR_Q0_1_INTRO_18_err_intro_q0_1_18;
assign err_intro_q0_1_frmC[19] =  o_LDPC_DEC_ERR_Q0_1_INTRO_19_err_intro_q0_1_19;
assign err_intro_q0_1_frmC[20] =  o_LDPC_DEC_ERR_Q0_1_INTRO_20_err_intro_q0_1_20;
assign err_intro_q0_1_frmC[21] =  o_LDPC_DEC_ERR_Q0_1_INTRO_21_err_intro_q0_1_21;
assign err_intro_q0_1_frmC[22] =  o_LDPC_DEC_ERR_Q0_1_INTRO_22_err_intro_q0_1_22;
assign err_intro_q0_1_frmC[23] =  o_LDPC_DEC_ERR_Q0_1_INTRO_23_err_intro_q0_1_23;
assign err_intro_q0_1_frmC[24] =  o_LDPC_DEC_ERR_Q0_1_INTRO_24_err_intro_q0_1_24;
assign err_intro_q0_1_frmC[25] =  o_LDPC_DEC_ERR_Q0_1_INTRO_25_err_intro_q0_1_25;
assign err_intro_q0_1_frmC[26] =  o_LDPC_DEC_ERR_Q0_1_INTRO_26_err_intro_q0_1_26;
assign err_intro_q0_1_frmC[27] =  o_LDPC_DEC_ERR_Q0_1_INTRO_27_err_intro_q0_1_27;
assign err_intro_q0_1_frmC[28] =  o_LDPC_DEC_ERR_Q0_1_INTRO_28_err_intro_q0_1_28;
assign err_intro_q0_1_frmC[29] =  o_LDPC_DEC_ERR_Q0_1_INTRO_29_err_intro_q0_1_29;
assign err_intro_q0_1_frmC[30] =  o_LDPC_DEC_ERR_Q0_1_INTRO_30_err_intro_q0_1_30;
assign err_intro_q0_1_frmC[31] =  o_LDPC_DEC_ERR_Q0_1_INTRO_31_err_intro_q0_1_31;
assign err_intro_q0_1_frmC[32] =  o_LDPC_DEC_ERR_Q0_1_INTRO_32_err_intro_q0_1_32;
assign err_intro_q0_1_frmC[33] =  o_LDPC_DEC_ERR_Q0_1_INTRO_33_err_intro_q0_1_33;
assign err_intro_q0_1_frmC[34] =  o_LDPC_DEC_ERR_Q0_1_INTRO_34_err_intro_q0_1_34;
assign err_intro_q0_1_frmC[35] =  o_LDPC_DEC_ERR_Q0_1_INTRO_35_err_intro_q0_1_35;
assign err_intro_q0_1_frmC[36] =  o_LDPC_DEC_ERR_Q0_1_INTRO_36_err_intro_q0_1_36;
assign err_intro_q0_1_frmC[37] =  o_LDPC_DEC_ERR_Q0_1_INTRO_37_err_intro_q0_1_37;
assign err_intro_q0_1_frmC[38] =  o_LDPC_DEC_ERR_Q0_1_INTRO_38_err_intro_q0_1_38;
assign err_intro_q0_1_frmC[39] =  o_LDPC_DEC_ERR_Q0_1_INTRO_39_err_intro_q0_1_39;
assign err_intro_q0_1_frmC[40] =  o_LDPC_DEC_ERR_Q0_1_INTRO_40_err_intro_q0_1_40;
assign err_intro_q0_1_frmC[41] =  o_LDPC_DEC_ERR_Q0_1_INTRO_41_err_intro_q0_1_41;
assign err_intro_q0_1_frmC[42] =  o_LDPC_DEC_ERR_Q0_1_INTRO_42_err_intro_q0_1_42;
assign err_intro_q0_1_frmC[43] =  o_LDPC_DEC_ERR_Q0_1_INTRO_43_err_intro_q0_1_43;
assign err_intro_q0_1_frmC[44] =  o_LDPC_DEC_ERR_Q0_1_INTRO_44_err_intro_q0_1_44;
assign err_intro_q0_1_frmC[45] =  o_LDPC_DEC_ERR_Q0_1_INTRO_45_err_intro_q0_1_45;
assign err_intro_q0_1_frmC[46] =  o_LDPC_DEC_ERR_Q0_1_INTRO_46_err_intro_q0_1_46;
assign err_intro_q0_1_frmC[47] =  o_LDPC_DEC_ERR_Q0_1_INTRO_47_err_intro_q0_1_47;
assign err_intro_q0_1_frmC[48] =  o_LDPC_DEC_ERR_Q0_1_INTRO_48_err_intro_q0_1_48;
assign err_intro_q0_1_frmC[49] =  o_LDPC_DEC_ERR_Q0_1_INTRO_49_err_intro_q0_1_49;
assign err_intro_q0_1_frmC[50] =  o_LDPC_DEC_ERR_Q0_1_INTRO_50_err_intro_q0_1_50;
assign err_intro_q0_1_frmC[51] =  o_LDPC_DEC_ERR_Q0_1_INTRO_51_err_intro_q0_1_51;
assign err_intro_q0_1_frmC[52] =  o_LDPC_DEC_ERR_Q0_1_INTRO_52_err_intro_q0_1_52;
assign err_intro_q0_1_frmC[53] =  o_LDPC_DEC_ERR_Q0_1_INTRO_53_err_intro_q0_1_53;
assign err_intro_q0_1_frmC[54] =  o_LDPC_DEC_ERR_Q0_1_INTRO_54_err_intro_q0_1_54;
assign err_intro_q0_1_frmC[55] =  o_LDPC_DEC_ERR_Q0_1_INTRO_55_err_intro_q0_1_55;
assign err_intro_q0_1_frmC[56] =  o_LDPC_DEC_ERR_Q0_1_INTRO_56_err_intro_q0_1_56;
assign err_intro_q0_1_frmC[57] =  o_LDPC_DEC_ERR_Q0_1_INTRO_57_err_intro_q0_1_57;
assign err_intro_q0_1_frmC[58] =  o_LDPC_DEC_ERR_Q0_1_INTRO_58_err_intro_q0_1_58;
assign err_intro_q0_1_frmC[59] =  o_LDPC_DEC_ERR_Q0_1_INTRO_59_err_intro_q0_1_59;
assign err_intro_q0_1_frmC[60] =  o_LDPC_DEC_ERR_Q0_1_INTRO_60_err_intro_q0_1_60;
assign err_intro_q0_1_frmC[61] =  o_LDPC_DEC_ERR_Q0_1_INTRO_61_err_intro_q0_1_61;
assign err_intro_q0_1_frmC[62] =  o_LDPC_DEC_ERR_Q0_1_INTRO_62_err_intro_q0_1_62;
assign err_intro_q0_1_frmC[63] =  o_LDPC_DEC_ERR_Q0_1_INTRO_63_err_intro_q0_1_63;
assign err_intro_q0_1_frmC[64] =  o_LDPC_DEC_ERR_Q0_1_INTRO_64_err_intro_q0_1_64;
assign err_intro_q0_1_frmC[65] =  o_LDPC_DEC_ERR_Q0_1_INTRO_65_err_intro_q0_1_65;
assign err_intro_q0_1_frmC[66] =  o_LDPC_DEC_ERR_Q0_1_INTRO_66_err_intro_q0_1_66;
assign err_intro_q0_1_frmC[67] =  o_LDPC_DEC_ERR_Q0_1_INTRO_67_err_intro_q0_1_67;
assign err_intro_q0_1_frmC[68] =  o_LDPC_DEC_ERR_Q0_1_INTRO_68_err_intro_q0_1_68;
assign err_intro_q0_1_frmC[69] =  o_LDPC_DEC_ERR_Q0_1_INTRO_69_err_intro_q0_1_69;
assign err_intro_q0_1_frmC[70] =  o_LDPC_DEC_ERR_Q0_1_INTRO_70_err_intro_q0_1_70;
assign err_intro_q0_1_frmC[71] =  o_LDPC_DEC_ERR_Q0_1_INTRO_71_err_intro_q0_1_71;
assign err_intro_q0_1_frmC[72] =  o_LDPC_DEC_ERR_Q0_1_INTRO_72_err_intro_q0_1_72;
assign err_intro_q0_1_frmC[73] =  o_LDPC_DEC_ERR_Q0_1_INTRO_73_err_intro_q0_1_73;
assign err_intro_q0_1_frmC[74] =  o_LDPC_DEC_ERR_Q0_1_INTRO_74_err_intro_q0_1_74;
assign err_intro_q0_1_frmC[75] =  o_LDPC_DEC_ERR_Q0_1_INTRO_75_err_intro_q0_1_75;
assign err_intro_q0_1_frmC[76] =  o_LDPC_DEC_ERR_Q0_1_INTRO_76_err_intro_q0_1_76;
assign err_intro_q0_1_frmC[77] =  o_LDPC_DEC_ERR_Q0_1_INTRO_77_err_intro_q0_1_77;
assign err_intro_q0_1_frmC[78] =  o_LDPC_DEC_ERR_Q0_1_INTRO_78_err_intro_q0_1_78;
assign err_intro_q0_1_frmC[79] =  o_LDPC_DEC_ERR_Q0_1_INTRO_79_err_intro_q0_1_79;
assign err_intro_q0_1_frmC[80] =  o_LDPC_DEC_ERR_Q0_1_INTRO_80_err_intro_q0_1_80;
assign err_intro_q0_1_frmC[81] =  o_LDPC_DEC_ERR_Q0_1_INTRO_81_err_intro_q0_1_81;
assign err_intro_q0_1_frmC[82] =  o_LDPC_DEC_ERR_Q0_1_INTRO_82_err_intro_q0_1_82;
assign err_intro_q0_1_frmC[83] =  o_LDPC_DEC_ERR_Q0_1_INTRO_83_err_intro_q0_1_83;
assign err_intro_q0_1_frmC[84] =  o_LDPC_DEC_ERR_Q0_1_INTRO_84_err_intro_q0_1_84;
assign err_intro_q0_1_frmC[85] =  o_LDPC_DEC_ERR_Q0_1_INTRO_85_err_intro_q0_1_85;
assign err_intro_q0_1_frmC[86] =  o_LDPC_DEC_ERR_Q0_1_INTRO_86_err_intro_q0_1_86;
assign err_intro_q0_1_frmC[87] =  o_LDPC_DEC_ERR_Q0_1_INTRO_87_err_intro_q0_1_87;
assign err_intro_q0_1_frmC[88] =  o_LDPC_DEC_ERR_Q0_1_INTRO_88_err_intro_q0_1_88;
assign err_intro_q0_1_frmC[89] =  o_LDPC_DEC_ERR_Q0_1_INTRO_89_err_intro_q0_1_89;
assign err_intro_q0_1_frmC[90] =  o_LDPC_DEC_ERR_Q0_1_INTRO_90_err_intro_q0_1_90;
assign err_intro_q0_1_frmC[91] =  o_LDPC_DEC_ERR_Q0_1_INTRO_91_err_intro_q0_1_91;
assign err_intro_q0_1_frmC[92] =  o_LDPC_DEC_ERR_Q0_1_INTRO_92_err_intro_q0_1_92;
assign err_intro_q0_1_frmC[93] =  o_LDPC_DEC_ERR_Q0_1_INTRO_93_err_intro_q0_1_93;
assign err_intro_q0_1_frmC[94] =  o_LDPC_DEC_ERR_Q0_1_INTRO_94_err_intro_q0_1_94;
assign err_intro_q0_1_frmC[95] =  o_LDPC_DEC_ERR_Q0_1_INTRO_95_err_intro_q0_1_95;
assign err_intro_q0_1_frmC[96] =  o_LDPC_DEC_ERR_Q0_1_INTRO_96_err_intro_q0_1_96;
assign err_intro_q0_1_frmC[97] =  o_LDPC_DEC_ERR_Q0_1_INTRO_97_err_intro_q0_1_97;
assign err_intro_q0_1_frmC[98] =  o_LDPC_DEC_ERR_Q0_1_INTRO_98_err_intro_q0_1_98;
assign err_intro_q0_1_frmC[99] =  o_LDPC_DEC_ERR_Q0_1_INTRO_99_err_intro_q0_1_99;
assign err_intro_q0_1_frmC[100] =  o_LDPC_DEC_ERR_Q0_1_INTRO_100_err_intro_q0_1_100;
assign err_intro_q0_1_frmC[101] =  o_LDPC_DEC_ERR_Q0_1_INTRO_101_err_intro_q0_1_101;
assign err_intro_q0_1_frmC[102] =  o_LDPC_DEC_ERR_Q0_1_INTRO_102_err_intro_q0_1_102;
assign err_intro_q0_1_frmC[103] =  o_LDPC_DEC_ERR_Q0_1_INTRO_103_err_intro_q0_1_103;
assign err_intro_q0_1_frmC[104] =  o_LDPC_DEC_ERR_Q0_1_INTRO_104_err_intro_q0_1_104;
assign err_intro_q0_1_frmC[105] =  o_LDPC_DEC_ERR_Q0_1_INTRO_105_err_intro_q0_1_105;
assign err_intro_q0_1_frmC[106] =  o_LDPC_DEC_ERR_Q0_1_INTRO_106_err_intro_q0_1_106;
assign err_intro_q0_1_frmC[107] =  o_LDPC_DEC_ERR_Q0_1_INTRO_107_err_intro_q0_1_107;
assign err_intro_q0_1_frmC[108] =  o_LDPC_DEC_ERR_Q0_1_INTRO_108_err_intro_q0_1_108;
assign err_intro_q0_1_frmC[109] =  o_LDPC_DEC_ERR_Q0_1_INTRO_109_err_intro_q0_1_109;
assign err_intro_q0_1_frmC[110] =  o_LDPC_DEC_ERR_Q0_1_INTRO_110_err_intro_q0_1_110;
assign err_intro_q0_1_frmC[111] =  o_LDPC_DEC_ERR_Q0_1_INTRO_111_err_intro_q0_1_111;
assign err_intro_q0_1_frmC[112] =  o_LDPC_DEC_ERR_Q0_1_INTRO_112_err_intro_q0_1_112;
assign err_intro_q0_1_frmC[113] =  o_LDPC_DEC_ERR_Q0_1_INTRO_113_err_intro_q0_1_113;
assign err_intro_q0_1_frmC[114] =  o_LDPC_DEC_ERR_Q0_1_INTRO_114_err_intro_q0_1_114;
assign err_intro_q0_1_frmC[115] =  o_LDPC_DEC_ERR_Q0_1_INTRO_115_err_intro_q0_1_115;
assign err_intro_q0_1_frmC[116] =  o_LDPC_DEC_ERR_Q0_1_INTRO_116_err_intro_q0_1_116;
assign err_intro_q0_1_frmC[117] =  o_LDPC_DEC_ERR_Q0_1_INTRO_117_err_intro_q0_1_117;
assign err_intro_q0_1_frmC[118] =  o_LDPC_DEC_ERR_Q0_1_INTRO_118_err_intro_q0_1_118;
assign err_intro_q0_1_frmC[119] =  o_LDPC_DEC_ERR_Q0_1_INTRO_119_err_intro_q0_1_119;
assign err_intro_q0_1_frmC[120] =  o_LDPC_DEC_ERR_Q0_1_INTRO_120_err_intro_q0_1_120;
assign err_intro_q0_1_frmC[121] =  o_LDPC_DEC_ERR_Q0_1_INTRO_121_err_intro_q0_1_121;
assign err_intro_q0_1_frmC[122] =  o_LDPC_DEC_ERR_Q0_1_INTRO_122_err_intro_q0_1_122;
assign err_intro_q0_1_frmC[123] =  o_LDPC_DEC_ERR_Q0_1_INTRO_123_err_intro_q0_1_123;
assign err_intro_q0_1_frmC[124] =  o_LDPC_DEC_ERR_Q0_1_INTRO_124_err_intro_q0_1_124;
assign err_intro_q0_1_frmC[125] =  o_LDPC_DEC_ERR_Q0_1_INTRO_125_err_intro_q0_1_125;
assign err_intro_q0_1_frmC[126] =  o_LDPC_DEC_ERR_Q0_1_INTRO_126_err_intro_q0_1_126;
assign err_intro_q0_1_frmC[127] =  o_LDPC_DEC_ERR_Q0_1_INTRO_127_err_intro_q0_1_127;
assign err_intro_q0_1_frmC[128] =  o_LDPC_DEC_ERR_Q0_1_INTRO_128_err_intro_q0_1_128;
assign err_intro_q0_1_frmC[129] =  o_LDPC_DEC_ERR_Q0_1_INTRO_129_err_intro_q0_1_129;
assign err_intro_q0_1_frmC[130] =  o_LDPC_DEC_ERR_Q0_1_INTRO_130_err_intro_q0_1_130;
assign err_intro_q0_1_frmC[131] =  o_LDPC_DEC_ERR_Q0_1_INTRO_131_err_intro_q0_1_131;
assign err_intro_q0_1_frmC[132] =  o_LDPC_DEC_ERR_Q0_1_INTRO_132_err_intro_q0_1_132;
assign err_intro_q0_1_frmC[133] =  o_LDPC_DEC_ERR_Q0_1_INTRO_133_err_intro_q0_1_133;
assign err_intro_q0_1_frmC[134] =  o_LDPC_DEC_ERR_Q0_1_INTRO_134_err_intro_q0_1_134;
assign err_intro_q0_1_frmC[135] =  o_LDPC_DEC_ERR_Q0_1_INTRO_135_err_intro_q0_1_135;
assign err_intro_q0_1_frmC[136] =  o_LDPC_DEC_ERR_Q0_1_INTRO_136_err_intro_q0_1_136;
assign err_intro_q0_1_frmC[137] =  o_LDPC_DEC_ERR_Q0_1_INTRO_137_err_intro_q0_1_137;
assign err_intro_q0_1_frmC[138] =  o_LDPC_DEC_ERR_Q0_1_INTRO_138_err_intro_q0_1_138;
assign err_intro_q0_1_frmC[139] =  o_LDPC_DEC_ERR_Q0_1_INTRO_139_err_intro_q0_1_139;
assign err_intro_q0_1_frmC[140] =  o_LDPC_DEC_ERR_Q0_1_INTRO_140_err_intro_q0_1_140;
assign err_intro_q0_1_frmC[141] =  o_LDPC_DEC_ERR_Q0_1_INTRO_141_err_intro_q0_1_141;
assign err_intro_q0_1_frmC[142] =  o_LDPC_DEC_ERR_Q0_1_INTRO_142_err_intro_q0_1_142;
assign err_intro_q0_1_frmC[143] =  o_LDPC_DEC_ERR_Q0_1_INTRO_143_err_intro_q0_1_143;
assign err_intro_q0_1_frmC[144] =  o_LDPC_DEC_ERR_Q0_1_INTRO_144_err_intro_q0_1_144;
assign err_intro_q0_1_frmC[145] =  o_LDPC_DEC_ERR_Q0_1_INTRO_145_err_intro_q0_1_145;
assign err_intro_q0_1_frmC[146] =  o_LDPC_DEC_ERR_Q0_1_INTRO_146_err_intro_q0_1_146;
assign err_intro_q0_1_frmC[147] =  o_LDPC_DEC_ERR_Q0_1_INTRO_147_err_intro_q0_1_147;
assign err_intro_q0_1_frmC[148] =  o_LDPC_DEC_ERR_Q0_1_INTRO_148_err_intro_q0_1_148;
assign err_intro_q0_1_frmC[149] =  o_LDPC_DEC_ERR_Q0_1_INTRO_149_err_intro_q0_1_149;
assign err_intro_q0_1_frmC[150] =  o_LDPC_DEC_ERR_Q0_1_INTRO_150_err_intro_q0_1_150;
assign err_intro_q0_1_frmC[151] =  o_LDPC_DEC_ERR_Q0_1_INTRO_151_err_intro_q0_1_151;
assign err_intro_q0_1_frmC[152] =  o_LDPC_DEC_ERR_Q0_1_INTRO_152_err_intro_q0_1_152;
assign err_intro_q0_1_frmC[153] =  o_LDPC_DEC_ERR_Q0_1_INTRO_153_err_intro_q0_1_153;
assign err_intro_q0_1_frmC[154] =  o_LDPC_DEC_ERR_Q0_1_INTRO_154_err_intro_q0_1_154;
assign err_intro_q0_1_frmC[155] =  o_LDPC_DEC_ERR_Q0_1_INTRO_155_err_intro_q0_1_155;
assign err_intro_q0_1_frmC[156] =  o_LDPC_DEC_ERR_Q0_1_INTRO_156_err_intro_q0_1_156;
assign err_intro_q0_1_frmC[157] =  o_LDPC_DEC_ERR_Q0_1_INTRO_157_err_intro_q0_1_157;
assign err_intro_q0_1_frmC[158] =  o_LDPC_DEC_ERR_Q0_1_INTRO_158_err_intro_q0_1_158;
assign err_intro_q0_1_frmC[159] =  o_LDPC_DEC_ERR_Q0_1_INTRO_159_err_intro_q0_1_159;
assign err_intro_q0_1_frmC[160] =  o_LDPC_DEC_ERR_Q0_1_INTRO_160_err_intro_q0_1_160;
assign err_intro_q0_1_frmC[161] =  o_LDPC_DEC_ERR_Q0_1_INTRO_161_err_intro_q0_1_161;
assign err_intro_q0_1_frmC[162] =  o_LDPC_DEC_ERR_Q0_1_INTRO_162_err_intro_q0_1_162;
assign err_intro_q0_1_frmC[163] =  o_LDPC_DEC_ERR_Q0_1_INTRO_163_err_intro_q0_1_163;
assign err_intro_q0_1_frmC[164] =  o_LDPC_DEC_ERR_Q0_1_INTRO_164_err_intro_q0_1_164;
assign err_intro_q0_1_frmC[165] =  o_LDPC_DEC_ERR_Q0_1_INTRO_165_err_intro_q0_1_165;
assign err_intro_q0_1_frmC[166] =  o_LDPC_DEC_ERR_Q0_1_INTRO_166_err_intro_q0_1_166;
assign err_intro_q0_1_frmC[167] =  o_LDPC_DEC_ERR_Q0_1_INTRO_167_err_intro_q0_1_167;
assign err_intro_q0_1_frmC[168] =  o_LDPC_DEC_ERR_Q0_1_INTRO_168_err_intro_q0_1_168;
assign err_intro_q0_1_frmC[169] =  o_LDPC_DEC_ERR_Q0_1_INTRO_169_err_intro_q0_1_169;
assign err_intro_q0_1_frmC[170] =  o_LDPC_DEC_ERR_Q0_1_INTRO_170_err_intro_q0_1_170;
assign err_intro_q0_1_frmC[171] =  o_LDPC_DEC_ERR_Q0_1_INTRO_171_err_intro_q0_1_171;
assign err_intro_q0_1_frmC[172] =  o_LDPC_DEC_ERR_Q0_1_INTRO_172_err_intro_q0_1_172;
assign err_intro_q0_1_frmC[173] =  o_LDPC_DEC_ERR_Q0_1_INTRO_173_err_intro_q0_1_173;
assign err_intro_q0_1_frmC[174] =  o_LDPC_DEC_ERR_Q0_1_INTRO_174_err_intro_q0_1_174;
assign err_intro_q0_1_frmC[175] =  o_LDPC_DEC_ERR_Q0_1_INTRO_175_err_intro_q0_1_175;
assign err_intro_q0_1_frmC[176] =  o_LDPC_DEC_ERR_Q0_1_INTRO_176_err_intro_q0_1_176;
assign err_intro_q0_1_frmC[177] =  o_LDPC_DEC_ERR_Q0_1_INTRO_177_err_intro_q0_1_177;
assign err_intro_q0_1_frmC[178] =  o_LDPC_DEC_ERR_Q0_1_INTRO_178_err_intro_q0_1_178;
assign err_intro_q0_1_frmC[179] =  o_LDPC_DEC_ERR_Q0_1_INTRO_179_err_intro_q0_1_179;
assign err_intro_q0_1_frmC[180] =  o_LDPC_DEC_ERR_Q0_1_INTRO_180_err_intro_q0_1_180;
assign err_intro_q0_1_frmC[181] =  o_LDPC_DEC_ERR_Q0_1_INTRO_181_err_intro_q0_1_181;
assign err_intro_q0_1_frmC[182] =  o_LDPC_DEC_ERR_Q0_1_INTRO_182_err_intro_q0_1_182;
assign err_intro_q0_1_frmC[183] =  o_LDPC_DEC_ERR_Q0_1_INTRO_183_err_intro_q0_1_183;
assign err_intro_q0_1_frmC[184] =  o_LDPC_DEC_ERR_Q0_1_INTRO_184_err_intro_q0_1_184;
assign err_intro_q0_1_frmC[185] =  o_LDPC_DEC_ERR_Q0_1_INTRO_185_err_intro_q0_1_185;
assign err_intro_q0_1_frmC[186] =  o_LDPC_DEC_ERR_Q0_1_INTRO_186_err_intro_q0_1_186;
assign err_intro_q0_1_frmC[187] =  o_LDPC_DEC_ERR_Q0_1_INTRO_187_err_intro_q0_1_187;
assign err_intro_q0_1_frmC[188] =  o_LDPC_DEC_ERR_Q0_1_INTRO_188_err_intro_q0_1_188;
assign err_intro_q0_1_frmC[189] =  o_LDPC_DEC_ERR_Q0_1_INTRO_189_err_intro_q0_1_189;
assign err_intro_q0_1_frmC[190] =  o_LDPC_DEC_ERR_Q0_1_INTRO_190_err_intro_q0_1_190;
assign err_intro_q0_1_frmC[191] =  o_LDPC_DEC_ERR_Q0_1_INTRO_191_err_intro_q0_1_191;
assign err_intro_q0_1_frmC[192] =  o_LDPC_DEC_ERR_Q0_1_INTRO_192_err_intro_q0_1_192;
assign err_intro_q0_1_frmC[193] =  o_LDPC_DEC_ERR_Q0_1_INTRO_193_err_intro_q0_1_193;
assign err_intro_q0_1_frmC[194] =  o_LDPC_DEC_ERR_Q0_1_INTRO_194_err_intro_q0_1_194;
assign err_intro_q0_1_frmC[195] =  o_LDPC_DEC_ERR_Q0_1_INTRO_195_err_intro_q0_1_195;
assign err_intro_q0_1_frmC[196] =  o_LDPC_DEC_ERR_Q0_1_INTRO_196_err_intro_q0_1_196;
assign err_intro_q0_1_frmC[197] =  o_LDPC_DEC_ERR_Q0_1_INTRO_197_err_intro_q0_1_197;
assign err_intro_q0_1_frmC[198] =  o_LDPC_DEC_ERR_Q0_1_INTRO_198_err_intro_q0_1_198;
assign err_intro_q0_1_frmC[199] =  o_LDPC_DEC_ERR_Q0_1_INTRO_199_err_intro_q0_1_199;
assign err_intro_q0_1_frmC[200] =  o_LDPC_DEC_ERR_Q0_1_INTRO_200_err_intro_q0_1_200;
assign err_intro_q0_1_frmC[201] =  o_LDPC_DEC_ERR_Q0_1_INTRO_201_err_intro_q0_1_201;
assign err_intro_q0_1_frmC[202] =  o_LDPC_DEC_ERR_Q0_1_INTRO_202_err_intro_q0_1_202;
assign err_intro_q0_1_frmC[203] =  o_LDPC_DEC_ERR_Q0_1_INTRO_203_err_intro_q0_1_203;
assign err_intro_q0_1_frmC[204] =  o_LDPC_DEC_ERR_Q0_1_INTRO_204_err_intro_q0_1_204;
assign err_intro_q0_1_frmC[205] =  o_LDPC_DEC_ERR_Q0_1_INTRO_205_err_intro_q0_1_205;
assign err_intro_q0_1_frmC[206] =  o_LDPC_DEC_ERR_Q0_1_INTRO_206_err_intro_q0_1_206;
assign err_intro_q0_1_frmC[207] =  o_LDPC_DEC_ERR_Q0_1_INTRO_207_err_intro_q0_1_207;
assign err_intro =  o_LDPC_DEC_ERR_INTRODUCED_err_intro;
assign q0_0_frmC[   0] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_0_cword_q0_0 ;
 assign q0_0_frmC[   1] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_1_cword_q0_0 ;
 assign q0_0_frmC[   2] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_2_cword_q0_0 ;
 assign q0_0_frmC[   3] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_3_cword_q0_0 ;
 assign q0_0_frmC[   4] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_4_cword_q0_0 ;
 assign q0_0_frmC[   5] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_5_cword_q0_0 ;
 assign q0_0_frmC[   6] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_6_cword_q0_0 ;
 assign q0_0_frmC[   7] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_7_cword_q0_0 ;
 assign q0_0_frmC[   8] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_8_cword_q0_0 ;
 assign q0_0_frmC[   9] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_9_cword_q0_0 ;
 assign q0_0_frmC[   10] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_10_cword_q0_0 ;
 assign q0_0_frmC[   11] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_11_cword_q0_0 ;
 assign q0_0_frmC[   12] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_12_cword_q0_0 ;
 assign q0_0_frmC[   13] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_13_cword_q0_0 ;
 assign q0_0_frmC[   14] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_14_cword_q0_0 ;
 assign q0_0_frmC[   15] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_15_cword_q0_0 ;
 assign q0_0_frmC[   16] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_16_cword_q0_0 ;
 assign q0_0_frmC[   17] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_17_cword_q0_0 ;
 assign q0_0_frmC[   18] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_18_cword_q0_0 ;
 assign q0_0_frmC[   19] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_19_cword_q0_0 ;
 assign q0_0_frmC[   20] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_20_cword_q0_0 ;
 assign q0_0_frmC[   21] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_21_cword_q0_0 ;
 assign q0_0_frmC[   22] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_22_cword_q0_0 ;
 assign q0_0_frmC[   23] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_23_cword_q0_0 ;
 assign q0_0_frmC[   24] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_24_cword_q0_0 ;
 assign q0_0_frmC[   25] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_25_cword_q0_0 ;
 assign q0_0_frmC[   26] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_26_cword_q0_0 ;
 assign q0_0_frmC[   27] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_27_cword_q0_0 ;
 assign q0_0_frmC[   28] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_28_cword_q0_0 ;
 assign q0_0_frmC[   29] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_29_cword_q0_0 ;
 assign q0_0_frmC[   30] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_30_cword_q0_0 ;
 assign q0_0_frmC[   31] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_31_cword_q0_0 ;
 assign q0_0_frmC[   32] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_32_cword_q0_0 ;
 assign q0_0_frmC[   33] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_33_cword_q0_0 ;
 assign q0_0_frmC[   34] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_34_cword_q0_0 ;
 assign q0_0_frmC[   35] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_35_cword_q0_0 ;
 assign q0_0_frmC[   36] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_36_cword_q0_0 ;
 assign q0_0_frmC[   37] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_37_cword_q0_0 ;
 assign q0_0_frmC[   38] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_38_cword_q0_0 ;
 assign q0_0_frmC[   39] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_39_cword_q0_0 ;
 assign q0_0_frmC[   40] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_40_cword_q0_0 ;
 assign q0_0_frmC[   41] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_41_cword_q0_0 ;
 assign q0_0_frmC[   42] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_42_cword_q0_0 ;
 assign q0_0_frmC[   43] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_43_cword_q0_0 ;
 assign q0_0_frmC[   44] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_44_cword_q0_0 ;
 assign q0_0_frmC[   45] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_45_cword_q0_0 ;
 assign q0_0_frmC[   46] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_46_cword_q0_0 ;
 assign q0_0_frmC[   47] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_47_cword_q0_0 ;
 assign q0_0_frmC[   48] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_48_cword_q0_0 ;
 assign q0_0_frmC[   49] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_49_cword_q0_0 ;
 assign q0_0_frmC[   50] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_50_cword_q0_0 ;
 assign q0_0_frmC[   51] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_51_cword_q0_0 ;
 assign q0_0_frmC[   52] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_52_cword_q0_0 ;
 assign q0_0_frmC[   53] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_53_cword_q0_0 ;
 assign q0_0_frmC[   54] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_54_cword_q0_0 ;
 assign q0_0_frmC[   55] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_55_cword_q0_0 ;
 assign q0_0_frmC[   56] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_56_cword_q0_0 ;
 assign q0_0_frmC[   57] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_57_cword_q0_0 ;
 assign q0_0_frmC[   58] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_58_cword_q0_0 ;
 assign q0_0_frmC[   59] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_59_cword_q0_0 ;
 assign q0_0_frmC[   60] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_60_cword_q0_0 ;
 assign q0_0_frmC[   61] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_61_cword_q0_0 ;
 assign q0_0_frmC[   62] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_62_cword_q0_0 ;
 assign q0_0_frmC[   63] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_63_cword_q0_0 ;
 assign q0_0_frmC[   64] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_64_cword_q0_0 ;
 assign q0_0_frmC[   65] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_65_cword_q0_0 ;
 assign q0_0_frmC[   66] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_66_cword_q0_0 ;
 assign q0_0_frmC[   67] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_67_cword_q0_0 ;
 assign q0_0_frmC[   68] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_68_cword_q0_0 ;
 assign q0_0_frmC[   69] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_69_cword_q0_0 ;
 assign q0_0_frmC[   70] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_70_cword_q0_0 ;
 assign q0_0_frmC[   71] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_71_cword_q0_0 ;
 assign q0_0_frmC[   72] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_72_cword_q0_0 ;
 assign q0_0_frmC[   73] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_73_cword_q0_0 ;
 assign q0_0_frmC[   74] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_74_cword_q0_0 ;
 assign q0_0_frmC[   75] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_75_cword_q0_0 ;
 assign q0_0_frmC[   76] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_76_cword_q0_0 ;
 assign q0_0_frmC[   77] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_77_cword_q0_0 ;
 assign q0_0_frmC[   78] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_78_cword_q0_0 ;
 assign q0_0_frmC[   79] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_79_cword_q0_0 ;
 assign q0_0_frmC[   80] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_80_cword_q0_0 ;
 assign q0_0_frmC[   81] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_81_cword_q0_0 ;
 assign q0_0_frmC[   82] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_82_cword_q0_0 ;
 assign q0_0_frmC[   83] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_83_cword_q0_0 ;
 assign q0_0_frmC[   84] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_84_cword_q0_0 ;
 assign q0_0_frmC[   85] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_85_cword_q0_0 ;
 assign q0_0_frmC[   86] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_86_cword_q0_0 ;
 assign q0_0_frmC[   87] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_87_cword_q0_0 ;
 assign q0_0_frmC[   88] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_88_cword_q0_0 ;
 assign q0_0_frmC[   89] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_89_cword_q0_0 ;
 assign q0_0_frmC[   90] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_90_cword_q0_0 ;
 assign q0_0_frmC[   91] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_91_cword_q0_0 ;
 assign q0_0_frmC[   92] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_92_cword_q0_0 ;
 assign q0_0_frmC[   93] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_93_cword_q0_0 ;
 assign q0_0_frmC[   94] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_94_cword_q0_0 ;
 assign q0_0_frmC[   95] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_95_cword_q0_0 ;
 assign q0_0_frmC[   96] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_96_cword_q0_0 ;
 assign q0_0_frmC[   97] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_97_cword_q0_0 ;
 assign q0_0_frmC[   98] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_98_cword_q0_0 ;
 assign q0_0_frmC[   99] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_99_cword_q0_0 ;
 assign q0_0_frmC[   100] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_100_cword_q0_0 ;
 assign q0_0_frmC[   101] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_101_cword_q0_0 ;
 assign q0_0_frmC[   102] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_102_cword_q0_0 ;
 assign q0_0_frmC[   103] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_103_cword_q0_0 ;
 assign q0_0_frmC[   104] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_104_cword_q0_0 ;
 assign q0_0_frmC[   105] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_105_cword_q0_0 ;
 assign q0_0_frmC[   106] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_106_cword_q0_0 ;
 assign q0_0_frmC[   107] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_107_cword_q0_0 ;
 assign q0_0_frmC[   108] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_108_cword_q0_0 ;
 assign q0_0_frmC[   109] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_109_cword_q0_0 ;
 assign q0_0_frmC[   110] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_110_cword_q0_0 ;
 assign q0_0_frmC[   111] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_111_cword_q0_0 ;
 assign q0_0_frmC[   112] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_112_cword_q0_0 ;
 assign q0_0_frmC[   113] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_113_cword_q0_0 ;
 assign q0_0_frmC[   114] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_114_cword_q0_0 ;
 assign q0_0_frmC[   115] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_115_cword_q0_0 ;
 assign q0_0_frmC[   116] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_116_cword_q0_0 ;
 assign q0_0_frmC[   117] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_117_cword_q0_0 ;
 assign q0_0_frmC[   118] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_118_cword_q0_0 ;
 assign q0_0_frmC[   119] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_119_cword_q0_0 ;
 assign q0_0_frmC[   120] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_120_cword_q0_0 ;
 assign q0_0_frmC[   121] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_121_cword_q0_0 ;
 assign q0_0_frmC[   122] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_122_cword_q0_0 ;
 assign q0_0_frmC[   123] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_123_cword_q0_0 ;
 assign q0_0_frmC[   124] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_124_cword_q0_0 ;
 assign q0_0_frmC[   125] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_125_cword_q0_0 ;
 assign q0_0_frmC[   126] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_126_cword_q0_0 ;
 assign q0_0_frmC[   127] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_127_cword_q0_0 ;
 assign q0_0_frmC[   128] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_128_cword_q0_0 ;
 assign q0_0_frmC[   129] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_129_cword_q0_0 ;
 assign q0_0_frmC[   130] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_130_cword_q0_0 ;
 assign q0_0_frmC[   131] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_131_cword_q0_0 ;
 assign q0_0_frmC[   132] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_132_cword_q0_0 ;
 assign q0_0_frmC[   133] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_133_cword_q0_0 ;
 assign q0_0_frmC[   134] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_134_cword_q0_0 ;
 assign q0_0_frmC[   135] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_135_cword_q0_0 ;
 assign q0_0_frmC[   136] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_136_cword_q0_0 ;
 assign q0_0_frmC[   137] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_137_cword_q0_0 ;
 assign q0_0_frmC[   138] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_138_cword_q0_0 ;
 assign q0_0_frmC[   139] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_139_cword_q0_0 ;
 assign q0_0_frmC[   140] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_140_cword_q0_0 ;
 assign q0_0_frmC[   141] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_141_cword_q0_0 ;
 assign q0_0_frmC[   142] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_142_cword_q0_0 ;
 assign q0_0_frmC[   143] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_143_cword_q0_0 ;
 assign q0_0_frmC[   144] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_144_cword_q0_0 ;
 assign q0_0_frmC[   145] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_145_cword_q0_0 ;
 assign q0_0_frmC[   146] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_146_cword_q0_0 ;
 assign q0_0_frmC[   147] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_147_cword_q0_0 ;
 assign q0_0_frmC[   148] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_148_cword_q0_0 ;
 assign q0_0_frmC[   149] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_149_cword_q0_0 ;
 assign q0_0_frmC[   150] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_150_cword_q0_0 ;
 assign q0_0_frmC[   151] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_151_cword_q0_0 ;
 assign q0_0_frmC[   152] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_152_cword_q0_0 ;
 assign q0_0_frmC[   153] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_153_cword_q0_0 ;
 assign q0_0_frmC[   154] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_154_cword_q0_0 ;
 assign q0_0_frmC[   155] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_155_cword_q0_0 ;
 assign q0_0_frmC[   156] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_156_cword_q0_0 ;
 assign q0_0_frmC[   157] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_157_cword_q0_0 ;
 assign q0_0_frmC[   158] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_158_cword_q0_0 ;
 assign q0_0_frmC[   159] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_159_cword_q0_0 ;
 assign q0_0_frmC[   160] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_160_cword_q0_0 ;
 assign q0_0_frmC[   161] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_161_cword_q0_0 ;
 assign q0_0_frmC[   162] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_162_cword_q0_0 ;
 assign q0_0_frmC[   163] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_163_cword_q0_0 ;
 assign q0_0_frmC[   164] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_164_cword_q0_0 ;
 assign q0_0_frmC[   165] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_165_cword_q0_0 ;
 assign q0_0_frmC[   166] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_166_cword_q0_0 ;
 assign q0_0_frmC[   167] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_167_cword_q0_0 ;
 assign q0_0_frmC[   168] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_168_cword_q0_0 ;
 assign q0_0_frmC[   169] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_169_cword_q0_0 ;
 assign q0_0_frmC[   170] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_170_cword_q0_0 ;
 assign q0_0_frmC[   171] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_171_cword_q0_0 ;
 assign q0_0_frmC[   172] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_172_cword_q0_0 ;
 assign q0_0_frmC[   173] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_173_cword_q0_0 ;
 assign q0_0_frmC[   174] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_174_cword_q0_0 ;
 assign q0_0_frmC[   175] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_175_cword_q0_0 ;
 assign q0_0_frmC[   176] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_176_cword_q0_0 ;
 assign q0_0_frmC[   177] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_177_cword_q0_0 ;
 assign q0_0_frmC[   178] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_178_cword_q0_0 ;
 assign q0_0_frmC[   179] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_179_cword_q0_0 ;
 assign q0_0_frmC[   180] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_180_cword_q0_0 ;
 assign q0_0_frmC[   181] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_181_cword_q0_0 ;
 assign q0_0_frmC[   182] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_182_cword_q0_0 ;
 assign q0_0_frmC[   183] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_183_cword_q0_0 ;
 assign q0_0_frmC[   184] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_184_cword_q0_0 ;
 assign q0_0_frmC[   185] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_185_cword_q0_0 ;
 assign q0_0_frmC[   186] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_186_cword_q0_0 ;
 assign q0_0_frmC[   187] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_187_cword_q0_0 ;
 assign q0_0_frmC[   188] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_188_cword_q0_0 ;
 assign q0_0_frmC[   189] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_189_cword_q0_0 ;
 assign q0_0_frmC[   190] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_190_cword_q0_0 ;
 assign q0_0_frmC[   191] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_191_cword_q0_0 ;
 assign q0_0_frmC[   192] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_192_cword_q0_0 ;
 assign q0_0_frmC[   193] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_193_cword_q0_0 ;
 assign q0_0_frmC[   194] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_194_cword_q0_0 ;
 assign q0_0_frmC[   195] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_195_cword_q0_0 ;
 assign q0_0_frmC[   196] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_196_cword_q0_0 ;
 assign q0_0_frmC[   197] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_197_cword_q0_0 ;
 assign q0_0_frmC[   198] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_198_cword_q0_0 ;
 assign q0_0_frmC[   199] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_199_cword_q0_0 ;
 assign q0_0_frmC[   200] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_200_cword_q0_0 ;
 assign q0_0_frmC[   201] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_201_cword_q0_0 ;
 assign q0_0_frmC[   202] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_202_cword_q0_0 ;
 assign q0_0_frmC[   203] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_203_cword_q0_0 ;
 assign q0_0_frmC[   204] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_204_cword_q0_0 ;
 assign q0_0_frmC[   205] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_205_cword_q0_0 ;
 assign q0_0_frmC[   206] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_206_cword_q0_0 ;
 assign q0_0_frmC[   207] =  o_LDPC_DEC_CODEWRD_IN_Q0_0_207_cword_q0_0 ;
  assign q0_1_frmC[   0] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_0_cword_q0_1 ;
     assign q0_1_frmC[   1] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_1_cword_q0_1 ;
     assign q0_1_frmC[   2] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_2_cword_q0_1 ;
     assign q0_1_frmC[   3] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_3_cword_q0_1 ;
     assign q0_1_frmC[   4] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_4_cword_q0_1 ;
     assign q0_1_frmC[   5] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_5_cword_q0_1 ;
     assign q0_1_frmC[   6] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_6_cword_q0_1 ;
     assign q0_1_frmC[   7] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_7_cword_q0_1 ;
     assign q0_1_frmC[   8] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_8_cword_q0_1 ;
     assign q0_1_frmC[   9] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_9_cword_q0_1 ;
     assign q0_1_frmC[   10] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_10_cword_q0_1 ;
     assign q0_1_frmC[   11] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_11_cword_q0_1 ;
     assign q0_1_frmC[   12] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_12_cword_q0_1 ;
     assign q0_1_frmC[   13] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_13_cword_q0_1 ;
     assign q0_1_frmC[   14] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_14_cword_q0_1 ;
     assign q0_1_frmC[   15] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_15_cword_q0_1 ;
     assign q0_1_frmC[   16] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_16_cword_q0_1 ;
     assign q0_1_frmC[   17] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_17_cword_q0_1 ;
     assign q0_1_frmC[   18] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_18_cword_q0_1 ;
     assign q0_1_frmC[   19] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_19_cword_q0_1 ;
     assign q0_1_frmC[   20] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_20_cword_q0_1 ;
     assign q0_1_frmC[   21] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_21_cword_q0_1 ;
     assign q0_1_frmC[   22] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_22_cword_q0_1 ;
     assign q0_1_frmC[   23] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_23_cword_q0_1 ;
     assign q0_1_frmC[   24] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_24_cword_q0_1 ;
     assign q0_1_frmC[   25] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_25_cword_q0_1 ;
     assign q0_1_frmC[   26] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_26_cword_q0_1 ;
     assign q0_1_frmC[   27] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_27_cword_q0_1 ;
     assign q0_1_frmC[   28] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_28_cword_q0_1 ;
     assign q0_1_frmC[   29] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_29_cword_q0_1 ;
     assign q0_1_frmC[   30] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_30_cword_q0_1 ;
     assign q0_1_frmC[   31] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_31_cword_q0_1 ;
     assign q0_1_frmC[   32] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_32_cword_q0_1 ;
     assign q0_1_frmC[   33] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_33_cword_q0_1 ;
     assign q0_1_frmC[   34] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_34_cword_q0_1 ;
     assign q0_1_frmC[   35] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_35_cword_q0_1 ;
     assign q0_1_frmC[   36] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_36_cword_q0_1 ;
     assign q0_1_frmC[   37] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_37_cword_q0_1 ;
     assign q0_1_frmC[   38] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_38_cword_q0_1 ;
     assign q0_1_frmC[   39] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_39_cword_q0_1 ;
     assign q0_1_frmC[   40] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_40_cword_q0_1 ;
     assign q0_1_frmC[   41] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_41_cword_q0_1 ;
     assign q0_1_frmC[   42] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_42_cword_q0_1 ;
     assign q0_1_frmC[   43] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_43_cword_q0_1 ;
     assign q0_1_frmC[   44] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_44_cword_q0_1 ;
     assign q0_1_frmC[   45] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_45_cword_q0_1 ;
     assign q0_1_frmC[   46] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_46_cword_q0_1 ;
     assign q0_1_frmC[   47] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_47_cword_q0_1 ;
     assign q0_1_frmC[   48] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_48_cword_q0_1 ;
     assign q0_1_frmC[   49] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_49_cword_q0_1 ;
     assign q0_1_frmC[   50] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_50_cword_q0_1 ;
     assign q0_1_frmC[   51] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_51_cword_q0_1 ;
     assign q0_1_frmC[   52] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_52_cword_q0_1 ;
     assign q0_1_frmC[   53] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_53_cword_q0_1 ;
     assign q0_1_frmC[   54] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_54_cword_q0_1 ;
     assign q0_1_frmC[   55] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_55_cword_q0_1 ;
     assign q0_1_frmC[   56] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_56_cword_q0_1 ;
     assign q0_1_frmC[   57] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_57_cword_q0_1 ;
     assign q0_1_frmC[   58] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_58_cword_q0_1 ;
     assign q0_1_frmC[   59] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_59_cword_q0_1 ;
     assign q0_1_frmC[   60] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_60_cword_q0_1 ;
     assign q0_1_frmC[   61] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_61_cword_q0_1 ;
     assign q0_1_frmC[   62] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_62_cword_q0_1 ;
     assign q0_1_frmC[   63] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_63_cword_q0_1 ;
     assign q0_1_frmC[   64] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_64_cword_q0_1 ;
     assign q0_1_frmC[   65] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_65_cword_q0_1 ;
     assign q0_1_frmC[   66] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_66_cword_q0_1 ;
     assign q0_1_frmC[   67] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_67_cword_q0_1 ;
     assign q0_1_frmC[   68] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_68_cword_q0_1 ;
     assign q0_1_frmC[   69] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_69_cword_q0_1 ;
     assign q0_1_frmC[   70] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_70_cword_q0_1 ;
     assign q0_1_frmC[   71] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_71_cword_q0_1 ;
     assign q0_1_frmC[   72] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_72_cword_q0_1 ;
     assign q0_1_frmC[   73] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_73_cword_q0_1 ;
     assign q0_1_frmC[   74] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_74_cword_q0_1 ;
     assign q0_1_frmC[   75] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_75_cword_q0_1 ;
     assign q0_1_frmC[   76] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_76_cword_q0_1 ;
     assign q0_1_frmC[   77] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_77_cword_q0_1 ;
     assign q0_1_frmC[   78] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_78_cword_q0_1 ;
     assign q0_1_frmC[   79] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_79_cword_q0_1 ;
     assign q0_1_frmC[   80] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_80_cword_q0_1 ;
     assign q0_1_frmC[   81] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_81_cword_q0_1 ;
     assign q0_1_frmC[   82] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_82_cword_q0_1 ;
     assign q0_1_frmC[   83] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_83_cword_q0_1 ;
     assign q0_1_frmC[   84] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_84_cword_q0_1 ;
     assign q0_1_frmC[   85] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_85_cword_q0_1 ;
     assign q0_1_frmC[   86] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_86_cword_q0_1 ;
     assign q0_1_frmC[   87] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_87_cword_q0_1 ;
     assign q0_1_frmC[   88] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_88_cword_q0_1 ;
     assign q0_1_frmC[   89] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_89_cword_q0_1 ;
     assign q0_1_frmC[   90] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_90_cword_q0_1 ;
     assign q0_1_frmC[   91] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_91_cword_q0_1 ;
     assign q0_1_frmC[   92] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_92_cword_q0_1 ;
     assign q0_1_frmC[   93] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_93_cword_q0_1 ;
     assign q0_1_frmC[   94] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_94_cword_q0_1 ;
     assign q0_1_frmC[   95] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_95_cword_q0_1 ;
     assign q0_1_frmC[   96] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_96_cword_q0_1 ;
     assign q0_1_frmC[   97] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_97_cword_q0_1 ;
     assign q0_1_frmC[   98] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_98_cword_q0_1 ;
     assign q0_1_frmC[   99] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_99_cword_q0_1 ;
     assign q0_1_frmC[   100] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_100_cword_q0_1 ;
     assign q0_1_frmC[   101] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_101_cword_q0_1 ;
     assign q0_1_frmC[   102] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_102_cword_q0_1 ;
     assign q0_1_frmC[   103] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_103_cword_q0_1 ;
     assign q0_1_frmC[   104] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_104_cword_q0_1 ;
     assign q0_1_frmC[   105] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_105_cword_q0_1 ;
     assign q0_1_frmC[   106] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_106_cword_q0_1 ;
     assign q0_1_frmC[   107] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_107_cword_q0_1 ;
     assign q0_1_frmC[   108] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_108_cword_q0_1 ;
     assign q0_1_frmC[   109] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_109_cword_q0_1 ;
     assign q0_1_frmC[   110] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_110_cword_q0_1 ;
     assign q0_1_frmC[   111] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_111_cword_q0_1 ;
     assign q0_1_frmC[   112] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_112_cword_q0_1 ;
     assign q0_1_frmC[   113] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_113_cword_q0_1 ;
     assign q0_1_frmC[   114] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_114_cword_q0_1 ;
     assign q0_1_frmC[   115] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_115_cword_q0_1 ;
     assign q0_1_frmC[   116] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_116_cword_q0_1 ;
     assign q0_1_frmC[   117] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_117_cword_q0_1 ;
     assign q0_1_frmC[   118] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_118_cword_q0_1 ;
     assign q0_1_frmC[   119] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_119_cword_q0_1 ;
     assign q0_1_frmC[   120] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_120_cword_q0_1 ;
     assign q0_1_frmC[   121] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_121_cword_q0_1 ;
     assign q0_1_frmC[   122] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_122_cword_q0_1 ;
     assign q0_1_frmC[   123] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_123_cword_q0_1 ;
     assign q0_1_frmC[   124] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_124_cword_q0_1 ;
     assign q0_1_frmC[   125] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_125_cword_q0_1 ;
     assign q0_1_frmC[   126] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_126_cword_q0_1 ;
     assign q0_1_frmC[   127] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_127_cword_q0_1 ;
     assign q0_1_frmC[   128] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_128_cword_q0_1 ;
     assign q0_1_frmC[   129] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_129_cword_q0_1 ;
     assign q0_1_frmC[   130] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_130_cword_q0_1 ;
     assign q0_1_frmC[   131] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_131_cword_q0_1 ;
     assign q0_1_frmC[   132] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_132_cword_q0_1 ;
     assign q0_1_frmC[   133] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_133_cword_q0_1 ;
     assign q0_1_frmC[   134] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_134_cword_q0_1 ;
     assign q0_1_frmC[   135] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_135_cword_q0_1 ;
     assign q0_1_frmC[   136] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_136_cword_q0_1 ;
     assign q0_1_frmC[   137] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_137_cword_q0_1 ;
     assign q0_1_frmC[   138] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_138_cword_q0_1 ;
     assign q0_1_frmC[   139] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_139_cword_q0_1 ;
     assign q0_1_frmC[   140] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_140_cword_q0_1 ;
     assign q0_1_frmC[   141] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_141_cword_q0_1 ;
     assign q0_1_frmC[   142] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_142_cword_q0_1 ;
     assign q0_1_frmC[   143] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_143_cword_q0_1 ;
     assign q0_1_frmC[   144] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_144_cword_q0_1 ;
     assign q0_1_frmC[   145] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_145_cword_q0_1 ;
     assign q0_1_frmC[   146] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_146_cword_q0_1 ;
     assign q0_1_frmC[   147] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_147_cword_q0_1 ;
     assign q0_1_frmC[   148] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_148_cword_q0_1 ;
     assign q0_1_frmC[   149] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_149_cword_q0_1 ;
     assign q0_1_frmC[   150] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_150_cword_q0_1 ;
     assign q0_1_frmC[   151] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_151_cword_q0_1 ;
     assign q0_1_frmC[   152] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_152_cword_q0_1 ;
     assign q0_1_frmC[   153] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_153_cword_q0_1 ;
     assign q0_1_frmC[   154] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_154_cword_q0_1 ;
     assign q0_1_frmC[   155] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_155_cword_q0_1 ;
     assign q0_1_frmC[   156] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_156_cword_q0_1 ;
     assign q0_1_frmC[   157] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_157_cword_q0_1 ;
     assign q0_1_frmC[   158] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_158_cword_q0_1 ;
     assign q0_1_frmC[   159] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_159_cword_q0_1 ;
     assign q0_1_frmC[   160] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_160_cword_q0_1 ;
     assign q0_1_frmC[   161] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_161_cword_q0_1 ;
     assign q0_1_frmC[   162] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_162_cword_q0_1 ;
     assign q0_1_frmC[   163] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_163_cword_q0_1 ;
     assign q0_1_frmC[   164] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_164_cword_q0_1 ;
     assign q0_1_frmC[   165] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_165_cword_q0_1 ;
     assign q0_1_frmC[   166] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_166_cword_q0_1 ;
     assign q0_1_frmC[   167] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_167_cword_q0_1 ;
     assign q0_1_frmC[   168] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_168_cword_q0_1 ;
     assign q0_1_frmC[   169] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_169_cword_q0_1 ;
     assign q0_1_frmC[   170] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_170_cword_q0_1 ;
     assign q0_1_frmC[   171] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_171_cword_q0_1 ;
     assign q0_1_frmC[   172] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_172_cword_q0_1 ;
     assign q0_1_frmC[   173] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_173_cword_q0_1 ;
     assign q0_1_frmC[   174] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_174_cword_q0_1 ;
     assign q0_1_frmC[   175] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_175_cword_q0_1 ;
     assign q0_1_frmC[   176] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_176_cword_q0_1 ;
     assign q0_1_frmC[   177] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_177_cword_q0_1 ;
     assign q0_1_frmC[   178] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_178_cword_q0_1 ;
     assign q0_1_frmC[   179] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_179_cword_q0_1 ;
     assign q0_1_frmC[   180] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_180_cword_q0_1 ;
     assign q0_1_frmC[   181] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_181_cword_q0_1 ;
     assign q0_1_frmC[   182] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_182_cword_q0_1 ;
     assign q0_1_frmC[   183] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_183_cword_q0_1 ;
     assign q0_1_frmC[   184] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_184_cword_q0_1 ;
     assign q0_1_frmC[   185] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_185_cword_q0_1 ;
     assign q0_1_frmC[   186] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_186_cword_q0_1 ;
     assign q0_1_frmC[   187] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_187_cword_q0_1 ;
     assign q0_1_frmC[   188] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_188_cword_q0_1 ;
     assign q0_1_frmC[   189] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_189_cword_q0_1 ;
     assign q0_1_frmC[   190] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_190_cword_q0_1 ;
     assign q0_1_frmC[   191] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_191_cword_q0_1 ;
     assign q0_1_frmC[   192] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_192_cword_q0_1 ;
     assign q0_1_frmC[   193] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_193_cword_q0_1 ;
     assign q0_1_frmC[   194] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_194_cword_q0_1 ;
     assign q0_1_frmC[   195] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_195_cword_q0_1 ;
     assign q0_1_frmC[   196] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_196_cword_q0_1 ;
     assign q0_1_frmC[   197] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_197_cword_q0_1 ;
     assign q0_1_frmC[   198] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_198_cword_q0_1 ;
     assign q0_1_frmC[   199] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_199_cword_q0_1 ;
     assign q0_1_frmC[   200] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_200_cword_q0_1 ;
     assign q0_1_frmC[   201] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_201_cword_q0_1 ;
     assign q0_1_frmC[   202] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_202_cword_q0_1 ;
     assign q0_1_frmC[   203] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_203_cword_q0_1 ;
     assign q0_1_frmC[   204] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_204_cword_q0_1 ;
     assign q0_1_frmC[   205] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_205_cword_q0_1 ;
     assign q0_1_frmC[   206] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_206_cword_q0_1 ;
     assign q0_1_frmC[   207] =  o_LDPC_DEC_CODEWRD_IN_Q0_1_207_cword_q0_1 ;
    assign i_LDPC_DEC_ERR_INTRO_DECODER_err_intro_decoder_bit = err_intro_decoder;
assign percent_probability_int =  o_LDPC_DEC_PROBABILITY_perc_probability;
assign HamDist_loop_max =  o_LDPC_DEC_HAMDIST_LOOP_MAX_HamDist_loop_max;
assign HamDist_loop_percentage =  o_LDPC_DEC_HAMDIST_LOOP_PERCENTAGE_HamDist_loop_percentage;
assign HamDist_iir1 =  o_LDPC_DEC_HAMDIST_IIR1_HamDist_iir1;
assign HamDist_iir2 =  o_LDPC_DEC_HAMDIST_IIR2_NOT_USED_HamDist_iir2;
assign HamDist_iir3 =  o_LDPC_DEC_HAMDIST_IIR3_NOT_USED_HamDist_iir3;
assign i_LDPC_DEC_SYN_VALID_CWORD_DEC_FINAL_syn_valid_cword_dec = syn_valid_cword_dec ;
assign start_dec =  o_LDPC_DEC_START_DEC_start_dec;
assign i_LDPC_DEC_CONVERGED_LOOPS_ENDED_converged_loops_ended = converged_loops_ended;
assign reg_mprj_slave =  o_reg_mprj_slave_reg_mprj_slave;
assign i_LDPC_DEC_CONVERGED_PASS_FAIL_converged_pass_fail = converged_pass_fail;
assign i_LDPC_DEC_CODEWRD_OUT_BIT_0_final_cword = final_y_nr_dec[0];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_1_final_cword = final_y_nr_dec[1];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_2_final_cword = final_y_nr_dec[2];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_3_final_cword = final_y_nr_dec[3];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_4_final_cword = final_y_nr_dec[4];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_5_final_cword = final_y_nr_dec[5];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_6_final_cword = final_y_nr_dec[6];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_7_final_cword = final_y_nr_dec[7];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_8_final_cword = final_y_nr_dec[8];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_9_final_cword = final_y_nr_dec[9];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_10_final_cword = final_y_nr_dec[10];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_11_final_cword = final_y_nr_dec[11];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_12_final_cword = final_y_nr_dec[12];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_13_final_cword = final_y_nr_dec[13];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_14_final_cword = final_y_nr_dec[14];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_15_final_cword = final_y_nr_dec[15];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_16_final_cword = final_y_nr_dec[16];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_17_final_cword = final_y_nr_dec[17];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_18_final_cword = final_y_nr_dec[18];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_19_final_cword = final_y_nr_dec[19];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_20_final_cword = final_y_nr_dec[20];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_21_final_cword = final_y_nr_dec[21];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_22_final_cword = final_y_nr_dec[22];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_23_final_cword = final_y_nr_dec[23];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_24_final_cword = final_y_nr_dec[24];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_25_final_cword = final_y_nr_dec[25];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_26_final_cword = final_y_nr_dec[26];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_27_final_cword = final_y_nr_dec[27];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_28_final_cword = final_y_nr_dec[28];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_29_final_cword = final_y_nr_dec[29];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_30_final_cword = final_y_nr_dec[30];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_31_final_cword = final_y_nr_dec[31];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_32_final_cword = final_y_nr_dec[32];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_33_final_cword = final_y_nr_dec[33];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_34_final_cword = final_y_nr_dec[34];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_35_final_cword = final_y_nr_dec[35];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_36_final_cword = final_y_nr_dec[36];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_37_final_cword = final_y_nr_dec[37];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_38_final_cword = final_y_nr_dec[38];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_39_final_cword = final_y_nr_dec[39];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_40_final_cword = final_y_nr_dec[40];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_41_final_cword = final_y_nr_dec[41];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_42_final_cword = final_y_nr_dec[42];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_43_final_cword = final_y_nr_dec[43];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_44_final_cword = final_y_nr_dec[44];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_45_final_cword = final_y_nr_dec[45];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_46_final_cword = final_y_nr_dec[46];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_47_final_cword = final_y_nr_dec[47];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_48_final_cword = final_y_nr_dec[48];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_49_final_cword = final_y_nr_dec[49];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_50_final_cword = final_y_nr_dec[50];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_51_final_cword = final_y_nr_dec[51];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_52_final_cword = final_y_nr_dec[52];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_53_final_cword = final_y_nr_dec[53];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_54_final_cword = final_y_nr_dec[54];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_55_final_cword = final_y_nr_dec[55];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_56_final_cword = final_y_nr_dec[56];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_57_final_cword = final_y_nr_dec[57];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_58_final_cword = final_y_nr_dec[58];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_59_final_cword = final_y_nr_dec[59];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_60_final_cword = final_y_nr_dec[60];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_61_final_cword = final_y_nr_dec[61];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_62_final_cword = final_y_nr_dec[62];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_63_final_cword = final_y_nr_dec[63];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_64_final_cword = final_y_nr_dec[64];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_65_final_cword = final_y_nr_dec[65];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_66_final_cword = final_y_nr_dec[66];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_67_final_cword = final_y_nr_dec[67];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_68_final_cword = final_y_nr_dec[68];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_69_final_cword = final_y_nr_dec[69];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_70_final_cword = final_y_nr_dec[70];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_71_final_cword = final_y_nr_dec[71];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_72_final_cword = final_y_nr_dec[72];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_73_final_cword = final_y_nr_dec[73];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_74_final_cword = final_y_nr_dec[74];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_75_final_cword = final_y_nr_dec[75];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_76_final_cword = final_y_nr_dec[76];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_77_final_cword = final_y_nr_dec[77];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_78_final_cword = final_y_nr_dec[78];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_79_final_cword = final_y_nr_dec[79];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_80_final_cword = final_y_nr_dec[80];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_81_final_cword = final_y_nr_dec[81];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_82_final_cword = final_y_nr_dec[82];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_83_final_cword = final_y_nr_dec[83];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_84_final_cword = final_y_nr_dec[84];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_85_final_cword = final_y_nr_dec[85];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_86_final_cword = final_y_nr_dec[86];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_87_final_cword = final_y_nr_dec[87];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_88_final_cword = final_y_nr_dec[88];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_89_final_cword = final_y_nr_dec[89];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_90_final_cword = final_y_nr_dec[90];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_91_final_cword = final_y_nr_dec[91];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_92_final_cword = final_y_nr_dec[92];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_93_final_cword = final_y_nr_dec[93];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_94_final_cword = final_y_nr_dec[94];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_95_final_cword = final_y_nr_dec[95];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_96_final_cword = final_y_nr_dec[96];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_97_final_cword = final_y_nr_dec[97];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_98_final_cword = final_y_nr_dec[98];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_99_final_cword = final_y_nr_dec[99];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_100_final_cword = final_y_nr_dec[100];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_101_final_cword = final_y_nr_dec[101];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_102_final_cword = final_y_nr_dec[102];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_103_final_cword = final_y_nr_dec[103];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_104_final_cword = final_y_nr_dec[104];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_105_final_cword = final_y_nr_dec[105];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_106_final_cword = final_y_nr_dec[106];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_107_final_cword = final_y_nr_dec[107];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_108_final_cword = final_y_nr_dec[108];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_109_final_cword = final_y_nr_dec[109];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_110_final_cword = final_y_nr_dec[110];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_111_final_cword = final_y_nr_dec[111];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_112_final_cword = final_y_nr_dec[112];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_113_final_cword = final_y_nr_dec[113];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_114_final_cword = final_y_nr_dec[114];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_115_final_cword = final_y_nr_dec[115];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_116_final_cword = final_y_nr_dec[116];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_117_final_cword = final_y_nr_dec[117];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_118_final_cword = final_y_nr_dec[118];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_119_final_cword = final_y_nr_dec[119];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_120_final_cword = final_y_nr_dec[120];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_121_final_cword = final_y_nr_dec[121];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_122_final_cword = final_y_nr_dec[122];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_123_final_cword = final_y_nr_dec[123];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_124_final_cword = final_y_nr_dec[124];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_125_final_cword = final_y_nr_dec[125];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_126_final_cword = final_y_nr_dec[126];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_127_final_cword = final_y_nr_dec[127];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_128_final_cword = final_y_nr_dec[128];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_129_final_cword = final_y_nr_dec[129];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_130_final_cword = final_y_nr_dec[130];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_131_final_cword = final_y_nr_dec[131];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_132_final_cword = final_y_nr_dec[132];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_133_final_cword = final_y_nr_dec[133];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_134_final_cword = final_y_nr_dec[134];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_135_final_cword = final_y_nr_dec[135];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_136_final_cword = final_y_nr_dec[136];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_137_final_cword = final_y_nr_dec[137];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_138_final_cword = final_y_nr_dec[138];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_139_final_cword = final_y_nr_dec[139];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_140_final_cword = final_y_nr_dec[140];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_141_final_cword = final_y_nr_dec[141];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_142_final_cword = final_y_nr_dec[142];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_143_final_cword = final_y_nr_dec[143];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_144_final_cword = final_y_nr_dec[144];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_145_final_cword = final_y_nr_dec[145];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_146_final_cword = final_y_nr_dec[146];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_147_final_cword = final_y_nr_dec[147];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_148_final_cword = final_y_nr_dec[148];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_149_final_cword = final_y_nr_dec[149];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_150_final_cword = final_y_nr_dec[150];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_151_final_cword = final_y_nr_dec[151];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_152_final_cword = final_y_nr_dec[152];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_153_final_cword = final_y_nr_dec[153];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_154_final_cword = final_y_nr_dec[154];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_155_final_cword = final_y_nr_dec[155];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_156_final_cword = final_y_nr_dec[156];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_157_final_cword = final_y_nr_dec[157];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_158_final_cword = final_y_nr_dec[158];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_159_final_cword = final_y_nr_dec[159];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_160_final_cword = final_y_nr_dec[160];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_161_final_cword = final_y_nr_dec[161];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_162_final_cword = final_y_nr_dec[162];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_163_final_cword = final_y_nr_dec[163];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_164_final_cword = final_y_nr_dec[164];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_165_final_cword = final_y_nr_dec[165];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_166_final_cword = final_y_nr_dec[166];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_167_final_cword = final_y_nr_dec[167];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_168_final_cword = final_y_nr_dec[168];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_169_final_cword = final_y_nr_dec[169];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_170_final_cword = final_y_nr_dec[170];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_171_final_cword = final_y_nr_dec[171];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_172_final_cword = final_y_nr_dec[172];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_173_final_cword = final_y_nr_dec[173];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_174_final_cword = final_y_nr_dec[174];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_175_final_cword = final_y_nr_dec[175];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_176_final_cword = final_y_nr_dec[176];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_177_final_cword = final_y_nr_dec[177];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_178_final_cword = final_y_nr_dec[178];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_179_final_cword = final_y_nr_dec[179];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_180_final_cword = final_y_nr_dec[180];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_181_final_cword = final_y_nr_dec[181];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_182_final_cword = final_y_nr_dec[182];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_183_final_cword = final_y_nr_dec[183];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_184_final_cword = final_y_nr_dec[184];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_185_final_cword = final_y_nr_dec[185];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_186_final_cword = final_y_nr_dec[186];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_187_final_cword = final_y_nr_dec[187];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_188_final_cword = final_y_nr_dec[188];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_189_final_cword = final_y_nr_dec[189];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_190_final_cword = final_y_nr_dec[190];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_191_final_cword = final_y_nr_dec[191];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_192_final_cword = final_y_nr_dec[192];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_193_final_cword = final_y_nr_dec[193];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_194_final_cword = final_y_nr_dec[194];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_195_final_cword = final_y_nr_dec[195];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_196_final_cword = final_y_nr_dec[196];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_197_final_cword = final_y_nr_dec[197];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_198_final_cword = final_y_nr_dec[198];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_199_final_cword = final_y_nr_dec[199];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_200_final_cword = final_y_nr_dec[200];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_201_final_cword = final_y_nr_dec[201];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_202_final_cword = final_y_nr_dec[202];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_203_final_cword = final_y_nr_dec[203];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_204_final_cword = final_y_nr_dec[204];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_205_final_cword = final_y_nr_dec[205];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_206_final_cword = final_y_nr_dec[206];
assign i_LDPC_DEC_CODEWRD_OUT_BIT_207_final_cword = final_y_nr_dec[207];
assign pass_fail =  o_LDPC_DEC_PASS_FAIL_pass_fail;
assign i_LDPC_DEC_TB_PASS_FAIL_DECODER_tb_pass_fail_decoder_bit = tb_pass_fail_decoder;
