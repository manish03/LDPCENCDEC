version https://git-lfs.github.com/spec/v1
oid sha256:19352c6ee0821b7cc72f4649fa07aca0563e431e27165259b9e01018834c3fde
size 58483811
