package LDPC_CSR_ral_pkg;
  import uvm_pkg::*;
  import rggen_ral_pkg::*;
  `include "uvm_macros.svh"
  `include "rggen_ral_macros.svh"
  class LDPC_ENC_MSG_IN_0_reg_model extends rggen_ral_reg;
    rand rggen_ral_field msg_in;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(msg_in, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_MSG_IN_1_reg_model extends rggen_ral_reg;
    rand rggen_ral_field msg_in;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(msg_in, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_MSG_IN_2_reg_model extends rggen_ral_reg;
    rand rggen_ral_field msg_in;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(msg_in, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_MSG_IN_3_reg_model extends rggen_ral_reg;
    rand rggen_ral_field msg_in;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(msg_in, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_MSG_IN_4_reg_model extends rggen_ral_reg;
    rand rggen_ral_field msg_in;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(msg_in, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_MSG_IN_5_reg_model extends rggen_ral_reg;
    rand rggen_ral_field msg_in;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(msg_in, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_MSG_IN_6_reg_model extends rggen_ral_reg;
    rand rggen_ral_field msg_in;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(msg_in, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_MSG_IN_7_reg_model extends rggen_ral_reg;
    rand rggen_ral_field msg_in;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(msg_in, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_MSG_IN_8_reg_model extends rggen_ral_reg;
    rand rggen_ral_field msg_in;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(msg_in, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_MSG_IN_9_reg_model extends rggen_ral_reg;
    rand rggen_ral_field msg_in;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(msg_in, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_MSG_IN_10_reg_model extends rggen_ral_reg;
    rand rggen_ral_field msg_in;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(msg_in, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_MSG_IN_11_reg_model extends rggen_ral_reg;
    rand rggen_ral_field msg_in;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(msg_in, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_MSG_IN_12_reg_model extends rggen_ral_reg;
    rand rggen_ral_field msg_in;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(msg_in, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_MSG_IN_13_reg_model extends rggen_ral_reg;
    rand rggen_ral_field msg_in;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(msg_in, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_MSG_IN_14_reg_model extends rggen_ral_reg;
    rand rggen_ral_field msg_in;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(msg_in, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_MSG_IN_15_reg_model extends rggen_ral_reg;
    rand rggen_ral_field msg_in;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(msg_in, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_MSG_IN_16_reg_model extends rggen_ral_reg;
    rand rggen_ral_field msg_in;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(msg_in, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_MSG_IN_17_reg_model extends rggen_ral_reg;
    rand rggen_ral_field msg_in;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(msg_in, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_MSG_IN_18_reg_model extends rggen_ral_reg;
    rand rggen_ral_field msg_in;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(msg_in, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_MSG_IN_19_reg_model extends rggen_ral_reg;
    rand rggen_ral_field msg_in;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(msg_in, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_MSG_IN_20_reg_model extends rggen_ral_reg;
    rand rggen_ral_field msg_in;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(msg_in, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_MSG_IN_21_reg_model extends rggen_ral_reg;
    rand rggen_ral_field msg_in;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(msg_in, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_MSG_IN_22_reg_model extends rggen_ral_reg;
    rand rggen_ral_field msg_in;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(msg_in, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_MSG_IN_23_reg_model extends rggen_ral_reg;
    rand rggen_ral_field msg_in;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(msg_in, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_MSG_IN_24_reg_model extends rggen_ral_reg;
    rand rggen_ral_field msg_in;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(msg_in, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_MSG_IN_25_reg_model extends rggen_ral_reg;
    rand rggen_ral_field msg_in;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(msg_in, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_MSG_IN_26_reg_model extends rggen_ral_reg;
    rand rggen_ral_field msg_in;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(msg_in, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_MSG_IN_27_reg_model extends rggen_ral_reg;
    rand rggen_ral_field msg_in;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(msg_in, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_MSG_IN_28_reg_model extends rggen_ral_reg;
    rand rggen_ral_field msg_in;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(msg_in, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_MSG_IN_29_reg_model extends rggen_ral_reg;
    rand rggen_ral_field msg_in;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(msg_in, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_MSG_IN_30_reg_model extends rggen_ral_reg;
    rand rggen_ral_field msg_in;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(msg_in, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_MSG_IN_31_reg_model extends rggen_ral_reg;
    rand rggen_ral_field msg_in;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(msg_in, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_MSG_IN_32_reg_model extends rggen_ral_reg;
    rand rggen_ral_field msg_in;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(msg_in, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_MSG_IN_33_reg_model extends rggen_ral_reg;
    rand rggen_ral_field msg_in;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(msg_in, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_MSG_IN_34_reg_model extends rggen_ral_reg;
    rand rggen_ral_field msg_in;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(msg_in, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_MSG_IN_35_reg_model extends rggen_ral_reg;
    rand rggen_ral_field msg_in;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(msg_in, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_MSG_IN_36_reg_model extends rggen_ral_reg;
    rand rggen_ral_field msg_in;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(msg_in, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_MSG_IN_37_reg_model extends rggen_ral_reg;
    rand rggen_ral_field msg_in;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(msg_in, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_MSG_IN_38_reg_model extends rggen_ral_reg;
    rand rggen_ral_field msg_in;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(msg_in, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_MSG_IN_39_reg_model extends rggen_ral_reg;
    rand rggen_ral_field msg_in;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(msg_in, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_0_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_1_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_2_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_3_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_4_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_5_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_6_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_7_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_8_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_9_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_10_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_11_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_12_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_13_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_14_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_15_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_16_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_17_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_18_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_19_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_20_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_21_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_22_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_23_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_24_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_25_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_26_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_27_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_28_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_29_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_30_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_31_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_32_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_33_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_34_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_35_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_36_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_37_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_38_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_39_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_40_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_41_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_42_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_43_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_44_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_45_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_46_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_47_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_48_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_49_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_50_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_51_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_52_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_53_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_54_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_55_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_56_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_57_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_58_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_59_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_60_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_61_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_62_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_63_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_64_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_65_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_66_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_67_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_68_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_69_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_70_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_71_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_72_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_73_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_74_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_75_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_76_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_77_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_78_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_79_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_80_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_81_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_82_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_83_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_84_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_85_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_86_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_87_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_88_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_89_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_90_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_91_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_92_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_93_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_94_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_95_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_96_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_97_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_98_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_99_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_100_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_101_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_102_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_103_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_104_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_105_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_106_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_107_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_108_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_109_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_110_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_111_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_112_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_113_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_114_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_115_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_116_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_117_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_118_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_119_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_120_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_121_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_122_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_123_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_124_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_125_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_126_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_127_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_128_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_129_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_130_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_131_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_132_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_133_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_134_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_135_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_136_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_137_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_138_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_139_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_140_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_141_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_142_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_143_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_144_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_145_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_146_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_147_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_148_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_149_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_150_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_151_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_152_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_153_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_154_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_155_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_156_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_157_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_158_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_159_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_160_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_161_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_162_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_163_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_164_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_165_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_166_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_167_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_168_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_169_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_170_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_171_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_172_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_173_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_174_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_175_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_176_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_177_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_178_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_179_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_180_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_181_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_182_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_183_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_184_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_185_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_186_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_187_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_188_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_189_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_190_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_191_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_192_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_193_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_194_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_195_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_196_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_197_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_198_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_199_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_200_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_201_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_202_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_203_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_204_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_205_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_206_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_OUT_207_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_ENC_CODEWRD_VLD_reg_model extends rggen_ral_reg;
    rand rggen_ral_field enc_codeword_valid;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(enc_codeword_valid, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_SEL_FRMC_reg_model extends rggen_ral_reg;
    rand rggen_ral_field sel_q0_frmC;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(sel_q0_frmC, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_0_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_1_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_2_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_2;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_2, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_3_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_3;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_3, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_4_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_4;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_4, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_5_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_5;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_5, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_6_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_6;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_6, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_7_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_7;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_7, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_8_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_8;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_8, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_9_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_9;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_9, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_10_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_10;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_10, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_11_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_11;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_11, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_12_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_12;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_12, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_13_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_13;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_13, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_14_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_14;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_14, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_15_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_15;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_15, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_16_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_16;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_16, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_17_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_17;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_17, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_18_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_18;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_18, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_19_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_19;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_19, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_20_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_20;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_20, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_21_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_21;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_21, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_22_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_22;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_22, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_23_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_23;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_23, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_24_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_24;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_24, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_25_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_25;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_25, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_26_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_26;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_26, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_27_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_27;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_27, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_28_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_28;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_28, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_29_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_29;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_29, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_30_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_30;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_30, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_31_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_31;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_31, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_32_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_32;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_32, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_33_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_33;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_33, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_34_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_34;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_34, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_35_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_35;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_35, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_36_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_36;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_36, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_37_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_37;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_37, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_38_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_38;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_38, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_39_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_39;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_39, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_40_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_40;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_40, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_41_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_41;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_41, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_42_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_42;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_42, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_43_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_43;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_43, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_44_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_44;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_44, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_45_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_45;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_45, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_46_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_46;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_46, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_47_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_47;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_47, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_48_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_48;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_48, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_49_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_49;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_49, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_50_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_50;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_50, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_51_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_51;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_51, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_52_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_52;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_52, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_53_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_53;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_53, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_54_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_54;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_54, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_55_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_55;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_55, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_56_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_56;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_56, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_57_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_57;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_57, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_58_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_58;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_58, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_59_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_59;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_59, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_60_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_60;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_60, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_61_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_61;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_61, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_62_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_62;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_62, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_63_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_63;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_63, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_64_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_64;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_64, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_65_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_65;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_65, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_66_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_66;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_66, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_67_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_67;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_67, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_68_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_68;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_68, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_69_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_69;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_69, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_70_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_70;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_70, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_71_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_71;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_71, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_72_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_72;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_72, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_73_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_73;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_73, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_74_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_74;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_74, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_75_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_75;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_75, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_76_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_76;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_76, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_77_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_77;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_77, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_78_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_78;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_78, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_79_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_79;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_79, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_80_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_80;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_80, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_81_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_81;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_81, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_82_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_82;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_82, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_83_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_83;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_83, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_84_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_84;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_84, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_85_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_85;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_85, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_86_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_86;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_86, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_87_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_87;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_87, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_88_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_88;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_88, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_89_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_89;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_89, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_90_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_90;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_90, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_91_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_91;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_91, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_92_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_92;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_92, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_93_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_93;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_93, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_94_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_94;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_94, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_95_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_95;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_95, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_96_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_96;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_96, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_97_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_97;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_97, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_98_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_98;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_98, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_99_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_99;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_99, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_100_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_100;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_100, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_101_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_101;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_101, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_102_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_102;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_102, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_103_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_103;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_103, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_104_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_104;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_104, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_105_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_105;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_105, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_106_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_106;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_106, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_107_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_107;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_107, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_108_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_108;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_108, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_109_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_109;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_109, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_110_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_110;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_110, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_111_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_111;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_111, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_112_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_112;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_112, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_113_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_113;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_113, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_114_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_114;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_114, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_115_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_115;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_115, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_116_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_116;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_116, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_117_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_117;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_117, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_118_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_118;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_118, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_119_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_119;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_119, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_120_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_120;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_120, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_121_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_121;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_121, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_122_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_122;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_122, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_123_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_123;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_123, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_124_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_124;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_124, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_125_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_125;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_125, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_126_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_126;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_126, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_127_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_127;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_127, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_128_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_128;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_128, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_129_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_129;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_129, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_130_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_130;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_130, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_131_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_131;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_131, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_132_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_132;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_132, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_133_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_133;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_133, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_134_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_134;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_134, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_135_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_135;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_135, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_136_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_136;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_136, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_137_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_137;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_137, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_138_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_138;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_138, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_139_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_139;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_139, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_140_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_140;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_140, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_141_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_141;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_141, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_142_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_142;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_142, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_143_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_143;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_143, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_144_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_144;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_144, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_145_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_145;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_145, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_146_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_146;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_146, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_147_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_147;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_147, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_148_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_148;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_148, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_149_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_149;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_149, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_150_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_150;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_150, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_151_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_151;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_151, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_152_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_152;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_152, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_153_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_153;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_153, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_154_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_154;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_154, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_155_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_155;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_155, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_156_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_156;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_156, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_157_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_157;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_157, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_158_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_158;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_158, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_159_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_159;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_159, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_160_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_160;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_160, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_161_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_161;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_161, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_162_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_162;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_162, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_163_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_163;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_163, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_164_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_164;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_164, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_165_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_165;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_165, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_166_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_166;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_166, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_167_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_167;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_167, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_168_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_168;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_168, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_169_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_169;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_169, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_170_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_170;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_170, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_171_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_171;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_171, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_172_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_172;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_172, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_173_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_173;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_173, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_174_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_174;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_174, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_175_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_175;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_175, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_176_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_176;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_176, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_177_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_177;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_177, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_178_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_178;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_178, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_179_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_179;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_179, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_180_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_180;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_180, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_181_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_181;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_181, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_182_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_182;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_182, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_183_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_183;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_183, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_184_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_184;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_184, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_185_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_185;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_185, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_186_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_186;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_186, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_187_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_187;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_187, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_188_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_188;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_188, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_189_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_189;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_189, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_190_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_190;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_190, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_191_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_191;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_191, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_192_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_192;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_192, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_193_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_193;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_193, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_194_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_194;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_194, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_195_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_195;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_195, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_196_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_196;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_196, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_197_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_197;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_197, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_198_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_198;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_198, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_199_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_199;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_199, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_200_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_200;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_200, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_201_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_201;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_201, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_202_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_202;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_202, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_203_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_203;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_203, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_204_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_204;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_204, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_205_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_205;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_205, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_206_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_206;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_206, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_0_INTRO_207_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_0_207;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_0_207, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_0_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_1_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_2_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_2;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_2, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_3_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_3;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_3, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_4_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_4;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_4, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_5_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_5;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_5, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_6_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_6;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_6, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_7_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_7;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_7, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_8_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_8;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_8, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_9_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_9;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_9, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_10_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_10;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_10, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_11_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_11;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_11, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_12_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_12;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_12, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_13_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_13;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_13, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_14_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_14;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_14, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_15_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_15;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_15, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_16_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_16;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_16, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_17_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_17;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_17, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_18_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_18;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_18, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_19_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_19;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_19, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_20_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_20;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_20, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_21_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_21;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_21, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_22_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_22;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_22, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_23_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_23;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_23, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_24_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_24;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_24, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_25_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_25;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_25, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_26_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_26;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_26, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_27_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_27;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_27, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_28_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_28;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_28, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_29_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_29;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_29, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_30_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_30;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_30, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_31_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_31;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_31, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_32_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_32;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_32, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_33_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_33;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_33, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_34_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_34;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_34, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_35_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_35;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_35, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_36_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_36;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_36, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_37_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_37;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_37, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_38_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_38;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_38, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_39_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_39;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_39, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_40_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_40;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_40, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_41_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_41;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_41, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_42_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_42;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_42, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_43_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_43;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_43, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_44_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_44;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_44, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_45_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_45;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_45, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_46_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_46;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_46, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_47_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_47;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_47, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_48_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_48;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_48, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_49_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_49;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_49, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_50_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_50;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_50, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_51_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_51;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_51, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_52_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_52;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_52, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_53_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_53;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_53, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_54_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_54;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_54, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_55_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_55;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_55, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_56_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_56;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_56, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_57_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_57;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_57, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_58_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_58;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_58, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_59_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_59;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_59, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_60_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_60;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_60, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_61_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_61;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_61, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_62_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_62;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_62, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_63_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_63;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_63, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_64_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_64;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_64, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_65_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_65;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_65, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_66_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_66;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_66, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_67_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_67;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_67, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_68_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_68;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_68, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_69_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_69;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_69, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_70_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_70;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_70, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_71_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_71;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_71, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_72_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_72;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_72, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_73_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_73;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_73, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_74_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_74;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_74, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_75_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_75;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_75, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_76_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_76;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_76, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_77_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_77;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_77, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_78_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_78;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_78, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_79_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_79;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_79, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_80_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_80;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_80, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_81_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_81;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_81, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_82_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_82;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_82, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_83_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_83;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_83, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_84_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_84;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_84, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_85_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_85;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_85, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_86_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_86;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_86, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_87_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_87;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_87, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_88_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_88;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_88, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_89_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_89;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_89, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_90_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_90;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_90, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_91_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_91;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_91, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_92_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_92;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_92, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_93_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_93;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_93, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_94_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_94;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_94, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_95_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_95;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_95, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_96_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_96;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_96, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_97_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_97;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_97, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_98_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_98;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_98, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_99_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_99;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_99, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_100_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_100;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_100, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_101_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_101;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_101, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_102_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_102;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_102, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_103_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_103;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_103, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_104_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_104;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_104, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_105_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_105;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_105, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_106_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_106;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_106, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_107_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_107;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_107, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_108_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_108;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_108, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_109_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_109;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_109, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_110_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_110;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_110, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_111_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_111;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_111, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_112_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_112;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_112, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_113_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_113;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_113, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_114_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_114;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_114, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_115_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_115;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_115, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_116_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_116;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_116, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_117_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_117;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_117, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_118_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_118;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_118, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_119_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_119;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_119, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_120_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_120;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_120, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_121_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_121;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_121, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_122_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_122;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_122, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_123_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_123;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_123, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_124_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_124;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_124, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_125_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_125;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_125, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_126_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_126;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_126, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_127_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_127;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_127, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_128_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_128;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_128, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_129_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_129;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_129, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_130_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_130;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_130, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_131_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_131;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_131, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_132_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_132;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_132, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_133_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_133;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_133, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_134_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_134;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_134, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_135_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_135;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_135, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_136_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_136;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_136, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_137_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_137;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_137, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_138_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_138;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_138, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_139_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_139;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_139, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_140_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_140;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_140, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_141_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_141;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_141, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_142_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_142;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_142, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_143_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_143;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_143, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_144_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_144;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_144, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_145_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_145;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_145, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_146_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_146;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_146, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_147_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_147;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_147, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_148_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_148;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_148, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_149_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_149;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_149, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_150_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_150;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_150, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_151_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_151;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_151, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_152_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_152;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_152, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_153_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_153;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_153, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_154_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_154;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_154, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_155_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_155;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_155, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_156_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_156;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_156, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_157_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_157;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_157, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_158_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_158;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_158, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_159_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_159;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_159, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_160_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_160;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_160, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_161_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_161;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_161, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_162_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_162;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_162, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_163_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_163;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_163, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_164_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_164;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_164, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_165_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_165;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_165, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_166_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_166;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_166, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_167_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_167;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_167, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_168_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_168;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_168, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_169_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_169;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_169, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_170_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_170;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_170, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_171_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_171;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_171, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_172_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_172;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_172, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_173_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_173;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_173, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_174_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_174;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_174, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_175_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_175;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_175, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_176_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_176;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_176, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_177_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_177;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_177, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_178_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_178;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_178, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_179_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_179;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_179, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_180_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_180;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_180, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_181_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_181;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_181, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_182_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_182;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_182, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_183_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_183;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_183, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_184_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_184;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_184, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_185_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_185;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_185, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_186_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_186;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_186, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_187_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_187;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_187, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_188_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_188;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_188, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_189_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_189;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_189, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_190_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_190;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_190, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_191_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_191;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_191, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_192_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_192;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_192, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_193_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_193;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_193, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_194_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_194;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_194, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_195_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_195;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_195, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_196_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_196;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_196, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_197_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_197;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_197, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_198_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_198;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_198, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_199_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_199;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_199, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_200_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_200;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_200, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_201_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_201;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_201, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_202_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_202;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_202, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_203_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_203;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_203, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_204_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_204;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_204, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_205_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_205;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_205, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_206_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_206;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_206, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_Q0_1_INTRO_207_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_q0_1_207;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_q0_1_207, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_ERR_INTRODUCED_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_0_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_1_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_2_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_3_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_4_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_5_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_6_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_7_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_8_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_9_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_10_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_11_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_12_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_13_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_14_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_15_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_16_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_17_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_18_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_19_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_20_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_21_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_22_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_23_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_24_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_25_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_26_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_27_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_28_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_29_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_30_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_31_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_32_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_33_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_34_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_35_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_36_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_37_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_38_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_39_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_40_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_41_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_42_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_43_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_44_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_45_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_46_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_47_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_48_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_49_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_50_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_51_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_52_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_53_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_54_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_55_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_56_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_57_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_58_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_59_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_60_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_61_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_62_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_63_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_64_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_65_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_66_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_67_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_68_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_69_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_70_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_71_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_72_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_73_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_74_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_75_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_76_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_77_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_78_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_79_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_80_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_81_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_82_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_83_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_84_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_85_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_86_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_87_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_88_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_89_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_90_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_91_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_92_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_93_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_94_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_95_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_96_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_97_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_98_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_99_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_100_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_101_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_102_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_103_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_104_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_105_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_106_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_107_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_108_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_109_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_110_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_111_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_112_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_113_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_114_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_115_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_116_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_117_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_118_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_119_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_120_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_121_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_122_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_123_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_124_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_125_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_126_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_127_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_128_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_129_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_130_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_131_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_132_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_133_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_134_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_135_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_136_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_137_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_138_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_139_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_140_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_141_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_142_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_143_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_144_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_145_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_146_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_147_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_148_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_149_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_150_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_151_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_152_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_153_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_154_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_155_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_156_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_157_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_158_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_159_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_160_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_161_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_162_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_163_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_164_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_165_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_166_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_167_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_168_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_169_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_170_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_171_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_172_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_173_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_174_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_175_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_176_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_177_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_178_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_179_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_180_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_181_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_182_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_183_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_184_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_185_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_186_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_187_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_188_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_189_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_190_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_191_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_192_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_193_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_194_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_195_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_196_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_197_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_198_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_199_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_200_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_201_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_202_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_203_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_204_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_205_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_206_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_0_207_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_0;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_0, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_0_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_1_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_2_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_3_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_4_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_5_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_6_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_7_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_8_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_9_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_10_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_11_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_12_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_13_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_14_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_15_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_16_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_17_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_18_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_19_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_20_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_21_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_22_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_23_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_24_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_25_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_26_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_27_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_28_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_29_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_30_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_31_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_32_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_33_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_34_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_35_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_36_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_37_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_38_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_39_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_40_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_41_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_42_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_43_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_44_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_45_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_46_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_47_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_48_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_49_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_50_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_51_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_52_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_53_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_54_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_55_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_56_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_57_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_58_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_59_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_60_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_61_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_62_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_63_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_64_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_65_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_66_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_67_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_68_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_69_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_70_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_71_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_72_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_73_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_74_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_75_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_76_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_77_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_78_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_79_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_80_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_81_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_82_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_83_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_84_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_85_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_86_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_87_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_88_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_89_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_90_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_91_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_92_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_93_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_94_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_95_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_96_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_97_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_98_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_99_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_100_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_101_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_102_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_103_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_104_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_105_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_106_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_107_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_108_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_109_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_110_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_111_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_112_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_113_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_114_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_115_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_116_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_117_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_118_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_119_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_120_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_121_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_122_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_123_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_124_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_125_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_126_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_127_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_128_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_129_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_130_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_131_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_132_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_133_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_134_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_135_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_136_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_137_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_138_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_139_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_140_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_141_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_142_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_143_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_144_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_145_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_146_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_147_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_148_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_149_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_150_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_151_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_152_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_153_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_154_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_155_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_156_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_157_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_158_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_159_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_160_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_161_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_162_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_163_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_164_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_165_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_166_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_167_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_168_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_169_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_170_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_171_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_172_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_173_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_174_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_175_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_176_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_177_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_178_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_179_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_180_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_181_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_182_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_183_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_184_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_185_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_186_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_187_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_188_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_189_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_190_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_191_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_192_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_193_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_194_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_195_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_196_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_197_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_198_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_199_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_200_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_201_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_202_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_203_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_204_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_205_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_206_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_IN_q0_1_207_reg_model extends rggen_ral_reg;
    rand rggen_ral_field cword_q0_1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(cword_q0_1, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_err_intro_decoder_reg_model extends rggen_ral_reg;
    rand rggen_ral_field err_intro_decoder_bit;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(err_intro_decoder_bit, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_0_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_1_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_2_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_3_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_4_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_5_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_6_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_7_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_8_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_9_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_10_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_11_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_12_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_13_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_14_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_15_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_16_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_17_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_18_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_19_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_20_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_21_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_22_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_23_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_24_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_25_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_26_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_27_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_28_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_29_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_30_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_31_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_32_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_33_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_34_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_35_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_36_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_37_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_38_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_39_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_40_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_41_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_42_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_43_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_44_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_45_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_46_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_47_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_48_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_49_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_50_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_51_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_52_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_53_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_54_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_55_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_56_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_57_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_58_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_59_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_60_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_61_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_62_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_63_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_64_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_65_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_66_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_67_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_68_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_69_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_70_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_71_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_72_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_73_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_74_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_75_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_76_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_77_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_78_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_79_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_80_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_81_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_82_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_83_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_84_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_85_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_86_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_87_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_88_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_89_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_90_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_91_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_92_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_93_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_94_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_95_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_96_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_97_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_98_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_99_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_100_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_101_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_102_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_103_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_104_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_105_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_106_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_107_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_108_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_109_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_110_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_111_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_112_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_113_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_114_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_115_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_116_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_117_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_118_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_119_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_120_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_121_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_122_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_123_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_124_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_125_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_126_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_127_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_128_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_129_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_130_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_131_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_132_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_133_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_134_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_135_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_136_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_137_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_138_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_139_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_140_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_141_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_142_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_143_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_144_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_145_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_146_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_147_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_148_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_149_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_150_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_151_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_152_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_153_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_154_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_155_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_156_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_157_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_158_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_159_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_160_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_161_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_162_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_163_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_164_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_165_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_166_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_EXPSYND_167_reg_model extends rggen_ral_reg;
    rand rggen_ral_field exp_syn;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(exp_syn, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_PROBABILITY_reg_model extends rggen_ral_reg;
    rand rggen_ral_field perc_probability;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(perc_probability, 0, 32, "RW", 0, 32'h00000000, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_HAMDIST_LOOP_MAX_reg_model extends rggen_ral_reg;
    rand rggen_ral_field HamDist_loop_max;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(HamDist_loop_max, 0, 32, "RW", 0, 32'h00000000, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_HAMDIST_LOOP_PERCENTAGE_reg_model extends rggen_ral_reg;
    rand rggen_ral_field HamDist_loop_percentage;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(HamDist_loop_percentage, 0, 32, "RW", 0, 32'h00000000, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_HAMDIST_IIR1_reg_model extends rggen_ral_reg;
    rand rggen_ral_field HamDist_iir1;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(HamDist_iir1, 0, 32, "RW", 0, 32'h00000000, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_HAMDIST_IIR2_NOT_USED_reg_model extends rggen_ral_reg;
    rand rggen_ral_field HamDist_iir2;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(HamDist_iir2, 0, 32, "RW", 0, 32'h00000000, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_HAMDIST_IIR3_NOT_USED_reg_model extends rggen_ral_reg;
    rand rggen_ral_field HamDist_iir3;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(HamDist_iir3, 0, 32, "RW", 0, 32'h00000000, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_SYN_VALID_CWORD_DEC_final_reg_model extends rggen_ral_reg;
    rand rggen_ral_field syn_valid_cword_dec;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(syn_valid_cword_dec, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_START_DEC_reg_model extends rggen_ral_reg;
    rand rggen_ral_field start_dec;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(start_dec, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CONVERGED_LOOPS_ENDED_reg_model extends rggen_ral_reg;
    rand rggen_ral_field converged_loops_ended;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(converged_loops_ended, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CONVERGED_PASS_FAIL_reg_model extends rggen_ral_reg;
    rand rggen_ral_field converged_pass_fail;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(converged_pass_fail, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_0_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_1_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_2_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_3_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_4_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_5_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_6_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_7_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_8_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_9_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_10_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_11_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_12_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_13_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_14_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_15_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_16_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_17_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_18_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_19_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_20_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_21_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_22_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_23_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_24_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_25_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_26_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_27_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_28_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_29_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_30_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_31_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_32_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_33_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_34_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_35_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_36_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_37_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_38_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_39_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_40_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_41_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_42_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_43_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_44_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_45_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_46_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_47_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_48_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_49_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_50_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_51_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_52_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_53_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_54_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_55_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_56_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_57_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_58_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_59_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_60_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_61_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_62_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_63_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_64_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_65_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_66_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_67_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_68_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_69_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_70_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_71_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_72_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_73_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_74_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_75_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_76_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_77_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_78_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_79_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_80_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_81_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_82_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_83_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_84_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_85_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_86_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_87_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_88_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_89_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_90_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_91_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_92_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_93_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_94_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_95_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_96_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_97_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_98_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_99_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_100_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_101_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_102_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_103_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_104_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_105_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_106_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_107_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_108_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_109_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_110_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_111_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_112_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_113_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_114_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_115_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_116_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_117_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_118_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_119_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_120_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_121_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_122_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_123_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_124_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_125_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_126_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_127_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_128_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_129_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_130_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_131_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_132_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_133_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_134_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_135_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_136_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_137_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_138_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_139_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_140_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_141_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_142_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_143_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_144_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_145_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_146_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_147_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_148_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_149_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_150_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_151_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_152_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_153_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_154_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_155_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_156_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_157_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_158_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_159_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_160_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_161_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_162_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_163_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_164_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_165_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_166_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_167_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_168_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_169_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_170_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_171_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_172_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_173_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_174_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_175_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_176_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_177_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_178_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_179_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_180_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_181_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_182_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_183_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_184_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_185_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_186_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_187_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_188_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_189_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_190_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_191_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_192_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_193_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_194_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_195_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_196_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_197_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_198_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_199_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_200_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_201_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_202_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_203_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_204_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_205_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_206_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_CODEWRD_OUT_BIT_207_reg_model extends rggen_ral_reg;
    rand rggen_ral_field final_cword;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(final_cword, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_PASS_FAIL_reg_model extends rggen_ral_reg;
    rand rggen_ral_field pass_fail;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(pass_fail, 0, 1, "RW", 0, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_DEC_pass_fail_decoder_reg_model extends rggen_ral_reg;
    rand rggen_ral_field pass_fail_decoder_bit;
    function new(string name);
      super.new(name, 32, 0);
    endfunction
    function void build();
      `rggen_ral_create_field(pass_fail_decoder_bit, 0, 1, "RO", 1, 1'h0, 1, -1, "")
    endfunction
  endclass
  class LDPC_CSR_block_model extends rggen_ral_block;
    rand LDPC_ENC_MSG_IN_0_reg_model LDPC_ENC_MSG_IN_0;
    rand LDPC_ENC_MSG_IN_1_reg_model LDPC_ENC_MSG_IN_1;
    rand LDPC_ENC_MSG_IN_2_reg_model LDPC_ENC_MSG_IN_2;
    rand LDPC_ENC_MSG_IN_3_reg_model LDPC_ENC_MSG_IN_3;
    rand LDPC_ENC_MSG_IN_4_reg_model LDPC_ENC_MSG_IN_4;
    rand LDPC_ENC_MSG_IN_5_reg_model LDPC_ENC_MSG_IN_5;
    rand LDPC_ENC_MSG_IN_6_reg_model LDPC_ENC_MSG_IN_6;
    rand LDPC_ENC_MSG_IN_7_reg_model LDPC_ENC_MSG_IN_7;
    rand LDPC_ENC_MSG_IN_8_reg_model LDPC_ENC_MSG_IN_8;
    rand LDPC_ENC_MSG_IN_9_reg_model LDPC_ENC_MSG_IN_9;
    rand LDPC_ENC_MSG_IN_10_reg_model LDPC_ENC_MSG_IN_10;
    rand LDPC_ENC_MSG_IN_11_reg_model LDPC_ENC_MSG_IN_11;
    rand LDPC_ENC_MSG_IN_12_reg_model LDPC_ENC_MSG_IN_12;
    rand LDPC_ENC_MSG_IN_13_reg_model LDPC_ENC_MSG_IN_13;
    rand LDPC_ENC_MSG_IN_14_reg_model LDPC_ENC_MSG_IN_14;
    rand LDPC_ENC_MSG_IN_15_reg_model LDPC_ENC_MSG_IN_15;
    rand LDPC_ENC_MSG_IN_16_reg_model LDPC_ENC_MSG_IN_16;
    rand LDPC_ENC_MSG_IN_17_reg_model LDPC_ENC_MSG_IN_17;
    rand LDPC_ENC_MSG_IN_18_reg_model LDPC_ENC_MSG_IN_18;
    rand LDPC_ENC_MSG_IN_19_reg_model LDPC_ENC_MSG_IN_19;
    rand LDPC_ENC_MSG_IN_20_reg_model LDPC_ENC_MSG_IN_20;
    rand LDPC_ENC_MSG_IN_21_reg_model LDPC_ENC_MSG_IN_21;
    rand LDPC_ENC_MSG_IN_22_reg_model LDPC_ENC_MSG_IN_22;
    rand LDPC_ENC_MSG_IN_23_reg_model LDPC_ENC_MSG_IN_23;
    rand LDPC_ENC_MSG_IN_24_reg_model LDPC_ENC_MSG_IN_24;
    rand LDPC_ENC_MSG_IN_25_reg_model LDPC_ENC_MSG_IN_25;
    rand LDPC_ENC_MSG_IN_26_reg_model LDPC_ENC_MSG_IN_26;
    rand LDPC_ENC_MSG_IN_27_reg_model LDPC_ENC_MSG_IN_27;
    rand LDPC_ENC_MSG_IN_28_reg_model LDPC_ENC_MSG_IN_28;
    rand LDPC_ENC_MSG_IN_29_reg_model LDPC_ENC_MSG_IN_29;
    rand LDPC_ENC_MSG_IN_30_reg_model LDPC_ENC_MSG_IN_30;
    rand LDPC_ENC_MSG_IN_31_reg_model LDPC_ENC_MSG_IN_31;
    rand LDPC_ENC_MSG_IN_32_reg_model LDPC_ENC_MSG_IN_32;
    rand LDPC_ENC_MSG_IN_33_reg_model LDPC_ENC_MSG_IN_33;
    rand LDPC_ENC_MSG_IN_34_reg_model LDPC_ENC_MSG_IN_34;
    rand LDPC_ENC_MSG_IN_35_reg_model LDPC_ENC_MSG_IN_35;
    rand LDPC_ENC_MSG_IN_36_reg_model LDPC_ENC_MSG_IN_36;
    rand LDPC_ENC_MSG_IN_37_reg_model LDPC_ENC_MSG_IN_37;
    rand LDPC_ENC_MSG_IN_38_reg_model LDPC_ENC_MSG_IN_38;
    rand LDPC_ENC_MSG_IN_39_reg_model LDPC_ENC_MSG_IN_39;
    rand LDPC_ENC_CODEWRD_OUT_0_reg_model LDPC_ENC_CODEWRD_OUT_0;
    rand LDPC_ENC_CODEWRD_OUT_1_reg_model LDPC_ENC_CODEWRD_OUT_1;
    rand LDPC_ENC_CODEWRD_OUT_2_reg_model LDPC_ENC_CODEWRD_OUT_2;
    rand LDPC_ENC_CODEWRD_OUT_3_reg_model LDPC_ENC_CODEWRD_OUT_3;
    rand LDPC_ENC_CODEWRD_OUT_4_reg_model LDPC_ENC_CODEWRD_OUT_4;
    rand LDPC_ENC_CODEWRD_OUT_5_reg_model LDPC_ENC_CODEWRD_OUT_5;
    rand LDPC_ENC_CODEWRD_OUT_6_reg_model LDPC_ENC_CODEWRD_OUT_6;
    rand LDPC_ENC_CODEWRD_OUT_7_reg_model LDPC_ENC_CODEWRD_OUT_7;
    rand LDPC_ENC_CODEWRD_OUT_8_reg_model LDPC_ENC_CODEWRD_OUT_8;
    rand LDPC_ENC_CODEWRD_OUT_9_reg_model LDPC_ENC_CODEWRD_OUT_9;
    rand LDPC_ENC_CODEWRD_OUT_10_reg_model LDPC_ENC_CODEWRD_OUT_10;
    rand LDPC_ENC_CODEWRD_OUT_11_reg_model LDPC_ENC_CODEWRD_OUT_11;
    rand LDPC_ENC_CODEWRD_OUT_12_reg_model LDPC_ENC_CODEWRD_OUT_12;
    rand LDPC_ENC_CODEWRD_OUT_13_reg_model LDPC_ENC_CODEWRD_OUT_13;
    rand LDPC_ENC_CODEWRD_OUT_14_reg_model LDPC_ENC_CODEWRD_OUT_14;
    rand LDPC_ENC_CODEWRD_OUT_15_reg_model LDPC_ENC_CODEWRD_OUT_15;
    rand LDPC_ENC_CODEWRD_OUT_16_reg_model LDPC_ENC_CODEWRD_OUT_16;
    rand LDPC_ENC_CODEWRD_OUT_17_reg_model LDPC_ENC_CODEWRD_OUT_17;
    rand LDPC_ENC_CODEWRD_OUT_18_reg_model LDPC_ENC_CODEWRD_OUT_18;
    rand LDPC_ENC_CODEWRD_OUT_19_reg_model LDPC_ENC_CODEWRD_OUT_19;
    rand LDPC_ENC_CODEWRD_OUT_20_reg_model LDPC_ENC_CODEWRD_OUT_20;
    rand LDPC_ENC_CODEWRD_OUT_21_reg_model LDPC_ENC_CODEWRD_OUT_21;
    rand LDPC_ENC_CODEWRD_OUT_22_reg_model LDPC_ENC_CODEWRD_OUT_22;
    rand LDPC_ENC_CODEWRD_OUT_23_reg_model LDPC_ENC_CODEWRD_OUT_23;
    rand LDPC_ENC_CODEWRD_OUT_24_reg_model LDPC_ENC_CODEWRD_OUT_24;
    rand LDPC_ENC_CODEWRD_OUT_25_reg_model LDPC_ENC_CODEWRD_OUT_25;
    rand LDPC_ENC_CODEWRD_OUT_26_reg_model LDPC_ENC_CODEWRD_OUT_26;
    rand LDPC_ENC_CODEWRD_OUT_27_reg_model LDPC_ENC_CODEWRD_OUT_27;
    rand LDPC_ENC_CODEWRD_OUT_28_reg_model LDPC_ENC_CODEWRD_OUT_28;
    rand LDPC_ENC_CODEWRD_OUT_29_reg_model LDPC_ENC_CODEWRD_OUT_29;
    rand LDPC_ENC_CODEWRD_OUT_30_reg_model LDPC_ENC_CODEWRD_OUT_30;
    rand LDPC_ENC_CODEWRD_OUT_31_reg_model LDPC_ENC_CODEWRD_OUT_31;
    rand LDPC_ENC_CODEWRD_OUT_32_reg_model LDPC_ENC_CODEWRD_OUT_32;
    rand LDPC_ENC_CODEWRD_OUT_33_reg_model LDPC_ENC_CODEWRD_OUT_33;
    rand LDPC_ENC_CODEWRD_OUT_34_reg_model LDPC_ENC_CODEWRD_OUT_34;
    rand LDPC_ENC_CODEWRD_OUT_35_reg_model LDPC_ENC_CODEWRD_OUT_35;
    rand LDPC_ENC_CODEWRD_OUT_36_reg_model LDPC_ENC_CODEWRD_OUT_36;
    rand LDPC_ENC_CODEWRD_OUT_37_reg_model LDPC_ENC_CODEWRD_OUT_37;
    rand LDPC_ENC_CODEWRD_OUT_38_reg_model LDPC_ENC_CODEWRD_OUT_38;
    rand LDPC_ENC_CODEWRD_OUT_39_reg_model LDPC_ENC_CODEWRD_OUT_39;
    rand LDPC_ENC_CODEWRD_OUT_40_reg_model LDPC_ENC_CODEWRD_OUT_40;
    rand LDPC_ENC_CODEWRD_OUT_41_reg_model LDPC_ENC_CODEWRD_OUT_41;
    rand LDPC_ENC_CODEWRD_OUT_42_reg_model LDPC_ENC_CODEWRD_OUT_42;
    rand LDPC_ENC_CODEWRD_OUT_43_reg_model LDPC_ENC_CODEWRD_OUT_43;
    rand LDPC_ENC_CODEWRD_OUT_44_reg_model LDPC_ENC_CODEWRD_OUT_44;
    rand LDPC_ENC_CODEWRD_OUT_45_reg_model LDPC_ENC_CODEWRD_OUT_45;
    rand LDPC_ENC_CODEWRD_OUT_46_reg_model LDPC_ENC_CODEWRD_OUT_46;
    rand LDPC_ENC_CODEWRD_OUT_47_reg_model LDPC_ENC_CODEWRD_OUT_47;
    rand LDPC_ENC_CODEWRD_OUT_48_reg_model LDPC_ENC_CODEWRD_OUT_48;
    rand LDPC_ENC_CODEWRD_OUT_49_reg_model LDPC_ENC_CODEWRD_OUT_49;
    rand LDPC_ENC_CODEWRD_OUT_50_reg_model LDPC_ENC_CODEWRD_OUT_50;
    rand LDPC_ENC_CODEWRD_OUT_51_reg_model LDPC_ENC_CODEWRD_OUT_51;
    rand LDPC_ENC_CODEWRD_OUT_52_reg_model LDPC_ENC_CODEWRD_OUT_52;
    rand LDPC_ENC_CODEWRD_OUT_53_reg_model LDPC_ENC_CODEWRD_OUT_53;
    rand LDPC_ENC_CODEWRD_OUT_54_reg_model LDPC_ENC_CODEWRD_OUT_54;
    rand LDPC_ENC_CODEWRD_OUT_55_reg_model LDPC_ENC_CODEWRD_OUT_55;
    rand LDPC_ENC_CODEWRD_OUT_56_reg_model LDPC_ENC_CODEWRD_OUT_56;
    rand LDPC_ENC_CODEWRD_OUT_57_reg_model LDPC_ENC_CODEWRD_OUT_57;
    rand LDPC_ENC_CODEWRD_OUT_58_reg_model LDPC_ENC_CODEWRD_OUT_58;
    rand LDPC_ENC_CODEWRD_OUT_59_reg_model LDPC_ENC_CODEWRD_OUT_59;
    rand LDPC_ENC_CODEWRD_OUT_60_reg_model LDPC_ENC_CODEWRD_OUT_60;
    rand LDPC_ENC_CODEWRD_OUT_61_reg_model LDPC_ENC_CODEWRD_OUT_61;
    rand LDPC_ENC_CODEWRD_OUT_62_reg_model LDPC_ENC_CODEWRD_OUT_62;
    rand LDPC_ENC_CODEWRD_OUT_63_reg_model LDPC_ENC_CODEWRD_OUT_63;
    rand LDPC_ENC_CODEWRD_OUT_64_reg_model LDPC_ENC_CODEWRD_OUT_64;
    rand LDPC_ENC_CODEWRD_OUT_65_reg_model LDPC_ENC_CODEWRD_OUT_65;
    rand LDPC_ENC_CODEWRD_OUT_66_reg_model LDPC_ENC_CODEWRD_OUT_66;
    rand LDPC_ENC_CODEWRD_OUT_67_reg_model LDPC_ENC_CODEWRD_OUT_67;
    rand LDPC_ENC_CODEWRD_OUT_68_reg_model LDPC_ENC_CODEWRD_OUT_68;
    rand LDPC_ENC_CODEWRD_OUT_69_reg_model LDPC_ENC_CODEWRD_OUT_69;
    rand LDPC_ENC_CODEWRD_OUT_70_reg_model LDPC_ENC_CODEWRD_OUT_70;
    rand LDPC_ENC_CODEWRD_OUT_71_reg_model LDPC_ENC_CODEWRD_OUT_71;
    rand LDPC_ENC_CODEWRD_OUT_72_reg_model LDPC_ENC_CODEWRD_OUT_72;
    rand LDPC_ENC_CODEWRD_OUT_73_reg_model LDPC_ENC_CODEWRD_OUT_73;
    rand LDPC_ENC_CODEWRD_OUT_74_reg_model LDPC_ENC_CODEWRD_OUT_74;
    rand LDPC_ENC_CODEWRD_OUT_75_reg_model LDPC_ENC_CODEWRD_OUT_75;
    rand LDPC_ENC_CODEWRD_OUT_76_reg_model LDPC_ENC_CODEWRD_OUT_76;
    rand LDPC_ENC_CODEWRD_OUT_77_reg_model LDPC_ENC_CODEWRD_OUT_77;
    rand LDPC_ENC_CODEWRD_OUT_78_reg_model LDPC_ENC_CODEWRD_OUT_78;
    rand LDPC_ENC_CODEWRD_OUT_79_reg_model LDPC_ENC_CODEWRD_OUT_79;
    rand LDPC_ENC_CODEWRD_OUT_80_reg_model LDPC_ENC_CODEWRD_OUT_80;
    rand LDPC_ENC_CODEWRD_OUT_81_reg_model LDPC_ENC_CODEWRD_OUT_81;
    rand LDPC_ENC_CODEWRD_OUT_82_reg_model LDPC_ENC_CODEWRD_OUT_82;
    rand LDPC_ENC_CODEWRD_OUT_83_reg_model LDPC_ENC_CODEWRD_OUT_83;
    rand LDPC_ENC_CODEWRD_OUT_84_reg_model LDPC_ENC_CODEWRD_OUT_84;
    rand LDPC_ENC_CODEWRD_OUT_85_reg_model LDPC_ENC_CODEWRD_OUT_85;
    rand LDPC_ENC_CODEWRD_OUT_86_reg_model LDPC_ENC_CODEWRD_OUT_86;
    rand LDPC_ENC_CODEWRD_OUT_87_reg_model LDPC_ENC_CODEWRD_OUT_87;
    rand LDPC_ENC_CODEWRD_OUT_88_reg_model LDPC_ENC_CODEWRD_OUT_88;
    rand LDPC_ENC_CODEWRD_OUT_89_reg_model LDPC_ENC_CODEWRD_OUT_89;
    rand LDPC_ENC_CODEWRD_OUT_90_reg_model LDPC_ENC_CODEWRD_OUT_90;
    rand LDPC_ENC_CODEWRD_OUT_91_reg_model LDPC_ENC_CODEWRD_OUT_91;
    rand LDPC_ENC_CODEWRD_OUT_92_reg_model LDPC_ENC_CODEWRD_OUT_92;
    rand LDPC_ENC_CODEWRD_OUT_93_reg_model LDPC_ENC_CODEWRD_OUT_93;
    rand LDPC_ENC_CODEWRD_OUT_94_reg_model LDPC_ENC_CODEWRD_OUT_94;
    rand LDPC_ENC_CODEWRD_OUT_95_reg_model LDPC_ENC_CODEWRD_OUT_95;
    rand LDPC_ENC_CODEWRD_OUT_96_reg_model LDPC_ENC_CODEWRD_OUT_96;
    rand LDPC_ENC_CODEWRD_OUT_97_reg_model LDPC_ENC_CODEWRD_OUT_97;
    rand LDPC_ENC_CODEWRD_OUT_98_reg_model LDPC_ENC_CODEWRD_OUT_98;
    rand LDPC_ENC_CODEWRD_OUT_99_reg_model LDPC_ENC_CODEWRD_OUT_99;
    rand LDPC_ENC_CODEWRD_OUT_100_reg_model LDPC_ENC_CODEWRD_OUT_100;
    rand LDPC_ENC_CODEWRD_OUT_101_reg_model LDPC_ENC_CODEWRD_OUT_101;
    rand LDPC_ENC_CODEWRD_OUT_102_reg_model LDPC_ENC_CODEWRD_OUT_102;
    rand LDPC_ENC_CODEWRD_OUT_103_reg_model LDPC_ENC_CODEWRD_OUT_103;
    rand LDPC_ENC_CODEWRD_OUT_104_reg_model LDPC_ENC_CODEWRD_OUT_104;
    rand LDPC_ENC_CODEWRD_OUT_105_reg_model LDPC_ENC_CODEWRD_OUT_105;
    rand LDPC_ENC_CODEWRD_OUT_106_reg_model LDPC_ENC_CODEWRD_OUT_106;
    rand LDPC_ENC_CODEWRD_OUT_107_reg_model LDPC_ENC_CODEWRD_OUT_107;
    rand LDPC_ENC_CODEWRD_OUT_108_reg_model LDPC_ENC_CODEWRD_OUT_108;
    rand LDPC_ENC_CODEWRD_OUT_109_reg_model LDPC_ENC_CODEWRD_OUT_109;
    rand LDPC_ENC_CODEWRD_OUT_110_reg_model LDPC_ENC_CODEWRD_OUT_110;
    rand LDPC_ENC_CODEWRD_OUT_111_reg_model LDPC_ENC_CODEWRD_OUT_111;
    rand LDPC_ENC_CODEWRD_OUT_112_reg_model LDPC_ENC_CODEWRD_OUT_112;
    rand LDPC_ENC_CODEWRD_OUT_113_reg_model LDPC_ENC_CODEWRD_OUT_113;
    rand LDPC_ENC_CODEWRD_OUT_114_reg_model LDPC_ENC_CODEWRD_OUT_114;
    rand LDPC_ENC_CODEWRD_OUT_115_reg_model LDPC_ENC_CODEWRD_OUT_115;
    rand LDPC_ENC_CODEWRD_OUT_116_reg_model LDPC_ENC_CODEWRD_OUT_116;
    rand LDPC_ENC_CODEWRD_OUT_117_reg_model LDPC_ENC_CODEWRD_OUT_117;
    rand LDPC_ENC_CODEWRD_OUT_118_reg_model LDPC_ENC_CODEWRD_OUT_118;
    rand LDPC_ENC_CODEWRD_OUT_119_reg_model LDPC_ENC_CODEWRD_OUT_119;
    rand LDPC_ENC_CODEWRD_OUT_120_reg_model LDPC_ENC_CODEWRD_OUT_120;
    rand LDPC_ENC_CODEWRD_OUT_121_reg_model LDPC_ENC_CODEWRD_OUT_121;
    rand LDPC_ENC_CODEWRD_OUT_122_reg_model LDPC_ENC_CODEWRD_OUT_122;
    rand LDPC_ENC_CODEWRD_OUT_123_reg_model LDPC_ENC_CODEWRD_OUT_123;
    rand LDPC_ENC_CODEWRD_OUT_124_reg_model LDPC_ENC_CODEWRD_OUT_124;
    rand LDPC_ENC_CODEWRD_OUT_125_reg_model LDPC_ENC_CODEWRD_OUT_125;
    rand LDPC_ENC_CODEWRD_OUT_126_reg_model LDPC_ENC_CODEWRD_OUT_126;
    rand LDPC_ENC_CODEWRD_OUT_127_reg_model LDPC_ENC_CODEWRD_OUT_127;
    rand LDPC_ENC_CODEWRD_OUT_128_reg_model LDPC_ENC_CODEWRD_OUT_128;
    rand LDPC_ENC_CODEWRD_OUT_129_reg_model LDPC_ENC_CODEWRD_OUT_129;
    rand LDPC_ENC_CODEWRD_OUT_130_reg_model LDPC_ENC_CODEWRD_OUT_130;
    rand LDPC_ENC_CODEWRD_OUT_131_reg_model LDPC_ENC_CODEWRD_OUT_131;
    rand LDPC_ENC_CODEWRD_OUT_132_reg_model LDPC_ENC_CODEWRD_OUT_132;
    rand LDPC_ENC_CODEWRD_OUT_133_reg_model LDPC_ENC_CODEWRD_OUT_133;
    rand LDPC_ENC_CODEWRD_OUT_134_reg_model LDPC_ENC_CODEWRD_OUT_134;
    rand LDPC_ENC_CODEWRD_OUT_135_reg_model LDPC_ENC_CODEWRD_OUT_135;
    rand LDPC_ENC_CODEWRD_OUT_136_reg_model LDPC_ENC_CODEWRD_OUT_136;
    rand LDPC_ENC_CODEWRD_OUT_137_reg_model LDPC_ENC_CODEWRD_OUT_137;
    rand LDPC_ENC_CODEWRD_OUT_138_reg_model LDPC_ENC_CODEWRD_OUT_138;
    rand LDPC_ENC_CODEWRD_OUT_139_reg_model LDPC_ENC_CODEWRD_OUT_139;
    rand LDPC_ENC_CODEWRD_OUT_140_reg_model LDPC_ENC_CODEWRD_OUT_140;
    rand LDPC_ENC_CODEWRD_OUT_141_reg_model LDPC_ENC_CODEWRD_OUT_141;
    rand LDPC_ENC_CODEWRD_OUT_142_reg_model LDPC_ENC_CODEWRD_OUT_142;
    rand LDPC_ENC_CODEWRD_OUT_143_reg_model LDPC_ENC_CODEWRD_OUT_143;
    rand LDPC_ENC_CODEWRD_OUT_144_reg_model LDPC_ENC_CODEWRD_OUT_144;
    rand LDPC_ENC_CODEWRD_OUT_145_reg_model LDPC_ENC_CODEWRD_OUT_145;
    rand LDPC_ENC_CODEWRD_OUT_146_reg_model LDPC_ENC_CODEWRD_OUT_146;
    rand LDPC_ENC_CODEWRD_OUT_147_reg_model LDPC_ENC_CODEWRD_OUT_147;
    rand LDPC_ENC_CODEWRD_OUT_148_reg_model LDPC_ENC_CODEWRD_OUT_148;
    rand LDPC_ENC_CODEWRD_OUT_149_reg_model LDPC_ENC_CODEWRD_OUT_149;
    rand LDPC_ENC_CODEWRD_OUT_150_reg_model LDPC_ENC_CODEWRD_OUT_150;
    rand LDPC_ENC_CODEWRD_OUT_151_reg_model LDPC_ENC_CODEWRD_OUT_151;
    rand LDPC_ENC_CODEWRD_OUT_152_reg_model LDPC_ENC_CODEWRD_OUT_152;
    rand LDPC_ENC_CODEWRD_OUT_153_reg_model LDPC_ENC_CODEWRD_OUT_153;
    rand LDPC_ENC_CODEWRD_OUT_154_reg_model LDPC_ENC_CODEWRD_OUT_154;
    rand LDPC_ENC_CODEWRD_OUT_155_reg_model LDPC_ENC_CODEWRD_OUT_155;
    rand LDPC_ENC_CODEWRD_OUT_156_reg_model LDPC_ENC_CODEWRD_OUT_156;
    rand LDPC_ENC_CODEWRD_OUT_157_reg_model LDPC_ENC_CODEWRD_OUT_157;
    rand LDPC_ENC_CODEWRD_OUT_158_reg_model LDPC_ENC_CODEWRD_OUT_158;
    rand LDPC_ENC_CODEWRD_OUT_159_reg_model LDPC_ENC_CODEWRD_OUT_159;
    rand LDPC_ENC_CODEWRD_OUT_160_reg_model LDPC_ENC_CODEWRD_OUT_160;
    rand LDPC_ENC_CODEWRD_OUT_161_reg_model LDPC_ENC_CODEWRD_OUT_161;
    rand LDPC_ENC_CODEWRD_OUT_162_reg_model LDPC_ENC_CODEWRD_OUT_162;
    rand LDPC_ENC_CODEWRD_OUT_163_reg_model LDPC_ENC_CODEWRD_OUT_163;
    rand LDPC_ENC_CODEWRD_OUT_164_reg_model LDPC_ENC_CODEWRD_OUT_164;
    rand LDPC_ENC_CODEWRD_OUT_165_reg_model LDPC_ENC_CODEWRD_OUT_165;
    rand LDPC_ENC_CODEWRD_OUT_166_reg_model LDPC_ENC_CODEWRD_OUT_166;
    rand LDPC_ENC_CODEWRD_OUT_167_reg_model LDPC_ENC_CODEWRD_OUT_167;
    rand LDPC_ENC_CODEWRD_OUT_168_reg_model LDPC_ENC_CODEWRD_OUT_168;
    rand LDPC_ENC_CODEWRD_OUT_169_reg_model LDPC_ENC_CODEWRD_OUT_169;
    rand LDPC_ENC_CODEWRD_OUT_170_reg_model LDPC_ENC_CODEWRD_OUT_170;
    rand LDPC_ENC_CODEWRD_OUT_171_reg_model LDPC_ENC_CODEWRD_OUT_171;
    rand LDPC_ENC_CODEWRD_OUT_172_reg_model LDPC_ENC_CODEWRD_OUT_172;
    rand LDPC_ENC_CODEWRD_OUT_173_reg_model LDPC_ENC_CODEWRD_OUT_173;
    rand LDPC_ENC_CODEWRD_OUT_174_reg_model LDPC_ENC_CODEWRD_OUT_174;
    rand LDPC_ENC_CODEWRD_OUT_175_reg_model LDPC_ENC_CODEWRD_OUT_175;
    rand LDPC_ENC_CODEWRD_OUT_176_reg_model LDPC_ENC_CODEWRD_OUT_176;
    rand LDPC_ENC_CODEWRD_OUT_177_reg_model LDPC_ENC_CODEWRD_OUT_177;
    rand LDPC_ENC_CODEWRD_OUT_178_reg_model LDPC_ENC_CODEWRD_OUT_178;
    rand LDPC_ENC_CODEWRD_OUT_179_reg_model LDPC_ENC_CODEWRD_OUT_179;
    rand LDPC_ENC_CODEWRD_OUT_180_reg_model LDPC_ENC_CODEWRD_OUT_180;
    rand LDPC_ENC_CODEWRD_OUT_181_reg_model LDPC_ENC_CODEWRD_OUT_181;
    rand LDPC_ENC_CODEWRD_OUT_182_reg_model LDPC_ENC_CODEWRD_OUT_182;
    rand LDPC_ENC_CODEWRD_OUT_183_reg_model LDPC_ENC_CODEWRD_OUT_183;
    rand LDPC_ENC_CODEWRD_OUT_184_reg_model LDPC_ENC_CODEWRD_OUT_184;
    rand LDPC_ENC_CODEWRD_OUT_185_reg_model LDPC_ENC_CODEWRD_OUT_185;
    rand LDPC_ENC_CODEWRD_OUT_186_reg_model LDPC_ENC_CODEWRD_OUT_186;
    rand LDPC_ENC_CODEWRD_OUT_187_reg_model LDPC_ENC_CODEWRD_OUT_187;
    rand LDPC_ENC_CODEWRD_OUT_188_reg_model LDPC_ENC_CODEWRD_OUT_188;
    rand LDPC_ENC_CODEWRD_OUT_189_reg_model LDPC_ENC_CODEWRD_OUT_189;
    rand LDPC_ENC_CODEWRD_OUT_190_reg_model LDPC_ENC_CODEWRD_OUT_190;
    rand LDPC_ENC_CODEWRD_OUT_191_reg_model LDPC_ENC_CODEWRD_OUT_191;
    rand LDPC_ENC_CODEWRD_OUT_192_reg_model LDPC_ENC_CODEWRD_OUT_192;
    rand LDPC_ENC_CODEWRD_OUT_193_reg_model LDPC_ENC_CODEWRD_OUT_193;
    rand LDPC_ENC_CODEWRD_OUT_194_reg_model LDPC_ENC_CODEWRD_OUT_194;
    rand LDPC_ENC_CODEWRD_OUT_195_reg_model LDPC_ENC_CODEWRD_OUT_195;
    rand LDPC_ENC_CODEWRD_OUT_196_reg_model LDPC_ENC_CODEWRD_OUT_196;
    rand LDPC_ENC_CODEWRD_OUT_197_reg_model LDPC_ENC_CODEWRD_OUT_197;
    rand LDPC_ENC_CODEWRD_OUT_198_reg_model LDPC_ENC_CODEWRD_OUT_198;
    rand LDPC_ENC_CODEWRD_OUT_199_reg_model LDPC_ENC_CODEWRD_OUT_199;
    rand LDPC_ENC_CODEWRD_OUT_200_reg_model LDPC_ENC_CODEWRD_OUT_200;
    rand LDPC_ENC_CODEWRD_OUT_201_reg_model LDPC_ENC_CODEWRD_OUT_201;
    rand LDPC_ENC_CODEWRD_OUT_202_reg_model LDPC_ENC_CODEWRD_OUT_202;
    rand LDPC_ENC_CODEWRD_OUT_203_reg_model LDPC_ENC_CODEWRD_OUT_203;
    rand LDPC_ENC_CODEWRD_OUT_204_reg_model LDPC_ENC_CODEWRD_OUT_204;
    rand LDPC_ENC_CODEWRD_OUT_205_reg_model LDPC_ENC_CODEWRD_OUT_205;
    rand LDPC_ENC_CODEWRD_OUT_206_reg_model LDPC_ENC_CODEWRD_OUT_206;
    rand LDPC_ENC_CODEWRD_OUT_207_reg_model LDPC_ENC_CODEWRD_OUT_207;
    rand LDPC_ENC_CODEWRD_VLD_reg_model LDPC_ENC_CODEWRD_VLD;
    rand LDPC_DEC_SEL_FRMC_reg_model LDPC_DEC_SEL_FRMC;
    rand LDPC_DEC_ERR_Q0_0_INTRO_0_reg_model LDPC_DEC_ERR_Q0_0_INTRO_0;
    rand LDPC_DEC_ERR_Q0_0_INTRO_1_reg_model LDPC_DEC_ERR_Q0_0_INTRO_1;
    rand LDPC_DEC_ERR_Q0_0_INTRO_2_reg_model LDPC_DEC_ERR_Q0_0_INTRO_2;
    rand LDPC_DEC_ERR_Q0_0_INTRO_3_reg_model LDPC_DEC_ERR_Q0_0_INTRO_3;
    rand LDPC_DEC_ERR_Q0_0_INTRO_4_reg_model LDPC_DEC_ERR_Q0_0_INTRO_4;
    rand LDPC_DEC_ERR_Q0_0_INTRO_5_reg_model LDPC_DEC_ERR_Q0_0_INTRO_5;
    rand LDPC_DEC_ERR_Q0_0_INTRO_6_reg_model LDPC_DEC_ERR_Q0_0_INTRO_6;
    rand LDPC_DEC_ERR_Q0_0_INTRO_7_reg_model LDPC_DEC_ERR_Q0_0_INTRO_7;
    rand LDPC_DEC_ERR_Q0_0_INTRO_8_reg_model LDPC_DEC_ERR_Q0_0_INTRO_8;
    rand LDPC_DEC_ERR_Q0_0_INTRO_9_reg_model LDPC_DEC_ERR_Q0_0_INTRO_9;
    rand LDPC_DEC_ERR_Q0_0_INTRO_10_reg_model LDPC_DEC_ERR_Q0_0_INTRO_10;
    rand LDPC_DEC_ERR_Q0_0_INTRO_11_reg_model LDPC_DEC_ERR_Q0_0_INTRO_11;
    rand LDPC_DEC_ERR_Q0_0_INTRO_12_reg_model LDPC_DEC_ERR_Q0_0_INTRO_12;
    rand LDPC_DEC_ERR_Q0_0_INTRO_13_reg_model LDPC_DEC_ERR_Q0_0_INTRO_13;
    rand LDPC_DEC_ERR_Q0_0_INTRO_14_reg_model LDPC_DEC_ERR_Q0_0_INTRO_14;
    rand LDPC_DEC_ERR_Q0_0_INTRO_15_reg_model LDPC_DEC_ERR_Q0_0_INTRO_15;
    rand LDPC_DEC_ERR_Q0_0_INTRO_16_reg_model LDPC_DEC_ERR_Q0_0_INTRO_16;
    rand LDPC_DEC_ERR_Q0_0_INTRO_17_reg_model LDPC_DEC_ERR_Q0_0_INTRO_17;
    rand LDPC_DEC_ERR_Q0_0_INTRO_18_reg_model LDPC_DEC_ERR_Q0_0_INTRO_18;
    rand LDPC_DEC_ERR_Q0_0_INTRO_19_reg_model LDPC_DEC_ERR_Q0_0_INTRO_19;
    rand LDPC_DEC_ERR_Q0_0_INTRO_20_reg_model LDPC_DEC_ERR_Q0_0_INTRO_20;
    rand LDPC_DEC_ERR_Q0_0_INTRO_21_reg_model LDPC_DEC_ERR_Q0_0_INTRO_21;
    rand LDPC_DEC_ERR_Q0_0_INTRO_22_reg_model LDPC_DEC_ERR_Q0_0_INTRO_22;
    rand LDPC_DEC_ERR_Q0_0_INTRO_23_reg_model LDPC_DEC_ERR_Q0_0_INTRO_23;
    rand LDPC_DEC_ERR_Q0_0_INTRO_24_reg_model LDPC_DEC_ERR_Q0_0_INTRO_24;
    rand LDPC_DEC_ERR_Q0_0_INTRO_25_reg_model LDPC_DEC_ERR_Q0_0_INTRO_25;
    rand LDPC_DEC_ERR_Q0_0_INTRO_26_reg_model LDPC_DEC_ERR_Q0_0_INTRO_26;
    rand LDPC_DEC_ERR_Q0_0_INTRO_27_reg_model LDPC_DEC_ERR_Q0_0_INTRO_27;
    rand LDPC_DEC_ERR_Q0_0_INTRO_28_reg_model LDPC_DEC_ERR_Q0_0_INTRO_28;
    rand LDPC_DEC_ERR_Q0_0_INTRO_29_reg_model LDPC_DEC_ERR_Q0_0_INTRO_29;
    rand LDPC_DEC_ERR_Q0_0_INTRO_30_reg_model LDPC_DEC_ERR_Q0_0_INTRO_30;
    rand LDPC_DEC_ERR_Q0_0_INTRO_31_reg_model LDPC_DEC_ERR_Q0_0_INTRO_31;
    rand LDPC_DEC_ERR_Q0_0_INTRO_32_reg_model LDPC_DEC_ERR_Q0_0_INTRO_32;
    rand LDPC_DEC_ERR_Q0_0_INTRO_33_reg_model LDPC_DEC_ERR_Q0_0_INTRO_33;
    rand LDPC_DEC_ERR_Q0_0_INTRO_34_reg_model LDPC_DEC_ERR_Q0_0_INTRO_34;
    rand LDPC_DEC_ERR_Q0_0_INTRO_35_reg_model LDPC_DEC_ERR_Q0_0_INTRO_35;
    rand LDPC_DEC_ERR_Q0_0_INTRO_36_reg_model LDPC_DEC_ERR_Q0_0_INTRO_36;
    rand LDPC_DEC_ERR_Q0_0_INTRO_37_reg_model LDPC_DEC_ERR_Q0_0_INTRO_37;
    rand LDPC_DEC_ERR_Q0_0_INTRO_38_reg_model LDPC_DEC_ERR_Q0_0_INTRO_38;
    rand LDPC_DEC_ERR_Q0_0_INTRO_39_reg_model LDPC_DEC_ERR_Q0_0_INTRO_39;
    rand LDPC_DEC_ERR_Q0_0_INTRO_40_reg_model LDPC_DEC_ERR_Q0_0_INTRO_40;
    rand LDPC_DEC_ERR_Q0_0_INTRO_41_reg_model LDPC_DEC_ERR_Q0_0_INTRO_41;
    rand LDPC_DEC_ERR_Q0_0_INTRO_42_reg_model LDPC_DEC_ERR_Q0_0_INTRO_42;
    rand LDPC_DEC_ERR_Q0_0_INTRO_43_reg_model LDPC_DEC_ERR_Q0_0_INTRO_43;
    rand LDPC_DEC_ERR_Q0_0_INTRO_44_reg_model LDPC_DEC_ERR_Q0_0_INTRO_44;
    rand LDPC_DEC_ERR_Q0_0_INTRO_45_reg_model LDPC_DEC_ERR_Q0_0_INTRO_45;
    rand LDPC_DEC_ERR_Q0_0_INTRO_46_reg_model LDPC_DEC_ERR_Q0_0_INTRO_46;
    rand LDPC_DEC_ERR_Q0_0_INTRO_47_reg_model LDPC_DEC_ERR_Q0_0_INTRO_47;
    rand LDPC_DEC_ERR_Q0_0_INTRO_48_reg_model LDPC_DEC_ERR_Q0_0_INTRO_48;
    rand LDPC_DEC_ERR_Q0_0_INTRO_49_reg_model LDPC_DEC_ERR_Q0_0_INTRO_49;
    rand LDPC_DEC_ERR_Q0_0_INTRO_50_reg_model LDPC_DEC_ERR_Q0_0_INTRO_50;
    rand LDPC_DEC_ERR_Q0_0_INTRO_51_reg_model LDPC_DEC_ERR_Q0_0_INTRO_51;
    rand LDPC_DEC_ERR_Q0_0_INTRO_52_reg_model LDPC_DEC_ERR_Q0_0_INTRO_52;
    rand LDPC_DEC_ERR_Q0_0_INTRO_53_reg_model LDPC_DEC_ERR_Q0_0_INTRO_53;
    rand LDPC_DEC_ERR_Q0_0_INTRO_54_reg_model LDPC_DEC_ERR_Q0_0_INTRO_54;
    rand LDPC_DEC_ERR_Q0_0_INTRO_55_reg_model LDPC_DEC_ERR_Q0_0_INTRO_55;
    rand LDPC_DEC_ERR_Q0_0_INTRO_56_reg_model LDPC_DEC_ERR_Q0_0_INTRO_56;
    rand LDPC_DEC_ERR_Q0_0_INTRO_57_reg_model LDPC_DEC_ERR_Q0_0_INTRO_57;
    rand LDPC_DEC_ERR_Q0_0_INTRO_58_reg_model LDPC_DEC_ERR_Q0_0_INTRO_58;
    rand LDPC_DEC_ERR_Q0_0_INTRO_59_reg_model LDPC_DEC_ERR_Q0_0_INTRO_59;
    rand LDPC_DEC_ERR_Q0_0_INTRO_60_reg_model LDPC_DEC_ERR_Q0_0_INTRO_60;
    rand LDPC_DEC_ERR_Q0_0_INTRO_61_reg_model LDPC_DEC_ERR_Q0_0_INTRO_61;
    rand LDPC_DEC_ERR_Q0_0_INTRO_62_reg_model LDPC_DEC_ERR_Q0_0_INTRO_62;
    rand LDPC_DEC_ERR_Q0_0_INTRO_63_reg_model LDPC_DEC_ERR_Q0_0_INTRO_63;
    rand LDPC_DEC_ERR_Q0_0_INTRO_64_reg_model LDPC_DEC_ERR_Q0_0_INTRO_64;
    rand LDPC_DEC_ERR_Q0_0_INTRO_65_reg_model LDPC_DEC_ERR_Q0_0_INTRO_65;
    rand LDPC_DEC_ERR_Q0_0_INTRO_66_reg_model LDPC_DEC_ERR_Q0_0_INTRO_66;
    rand LDPC_DEC_ERR_Q0_0_INTRO_67_reg_model LDPC_DEC_ERR_Q0_0_INTRO_67;
    rand LDPC_DEC_ERR_Q0_0_INTRO_68_reg_model LDPC_DEC_ERR_Q0_0_INTRO_68;
    rand LDPC_DEC_ERR_Q0_0_INTRO_69_reg_model LDPC_DEC_ERR_Q0_0_INTRO_69;
    rand LDPC_DEC_ERR_Q0_0_INTRO_70_reg_model LDPC_DEC_ERR_Q0_0_INTRO_70;
    rand LDPC_DEC_ERR_Q0_0_INTRO_71_reg_model LDPC_DEC_ERR_Q0_0_INTRO_71;
    rand LDPC_DEC_ERR_Q0_0_INTRO_72_reg_model LDPC_DEC_ERR_Q0_0_INTRO_72;
    rand LDPC_DEC_ERR_Q0_0_INTRO_73_reg_model LDPC_DEC_ERR_Q0_0_INTRO_73;
    rand LDPC_DEC_ERR_Q0_0_INTRO_74_reg_model LDPC_DEC_ERR_Q0_0_INTRO_74;
    rand LDPC_DEC_ERR_Q0_0_INTRO_75_reg_model LDPC_DEC_ERR_Q0_0_INTRO_75;
    rand LDPC_DEC_ERR_Q0_0_INTRO_76_reg_model LDPC_DEC_ERR_Q0_0_INTRO_76;
    rand LDPC_DEC_ERR_Q0_0_INTRO_77_reg_model LDPC_DEC_ERR_Q0_0_INTRO_77;
    rand LDPC_DEC_ERR_Q0_0_INTRO_78_reg_model LDPC_DEC_ERR_Q0_0_INTRO_78;
    rand LDPC_DEC_ERR_Q0_0_INTRO_79_reg_model LDPC_DEC_ERR_Q0_0_INTRO_79;
    rand LDPC_DEC_ERR_Q0_0_INTRO_80_reg_model LDPC_DEC_ERR_Q0_0_INTRO_80;
    rand LDPC_DEC_ERR_Q0_0_INTRO_81_reg_model LDPC_DEC_ERR_Q0_0_INTRO_81;
    rand LDPC_DEC_ERR_Q0_0_INTRO_82_reg_model LDPC_DEC_ERR_Q0_0_INTRO_82;
    rand LDPC_DEC_ERR_Q0_0_INTRO_83_reg_model LDPC_DEC_ERR_Q0_0_INTRO_83;
    rand LDPC_DEC_ERR_Q0_0_INTRO_84_reg_model LDPC_DEC_ERR_Q0_0_INTRO_84;
    rand LDPC_DEC_ERR_Q0_0_INTRO_85_reg_model LDPC_DEC_ERR_Q0_0_INTRO_85;
    rand LDPC_DEC_ERR_Q0_0_INTRO_86_reg_model LDPC_DEC_ERR_Q0_0_INTRO_86;
    rand LDPC_DEC_ERR_Q0_0_INTRO_87_reg_model LDPC_DEC_ERR_Q0_0_INTRO_87;
    rand LDPC_DEC_ERR_Q0_0_INTRO_88_reg_model LDPC_DEC_ERR_Q0_0_INTRO_88;
    rand LDPC_DEC_ERR_Q0_0_INTRO_89_reg_model LDPC_DEC_ERR_Q0_0_INTRO_89;
    rand LDPC_DEC_ERR_Q0_0_INTRO_90_reg_model LDPC_DEC_ERR_Q0_0_INTRO_90;
    rand LDPC_DEC_ERR_Q0_0_INTRO_91_reg_model LDPC_DEC_ERR_Q0_0_INTRO_91;
    rand LDPC_DEC_ERR_Q0_0_INTRO_92_reg_model LDPC_DEC_ERR_Q0_0_INTRO_92;
    rand LDPC_DEC_ERR_Q0_0_INTRO_93_reg_model LDPC_DEC_ERR_Q0_0_INTRO_93;
    rand LDPC_DEC_ERR_Q0_0_INTRO_94_reg_model LDPC_DEC_ERR_Q0_0_INTRO_94;
    rand LDPC_DEC_ERR_Q0_0_INTRO_95_reg_model LDPC_DEC_ERR_Q0_0_INTRO_95;
    rand LDPC_DEC_ERR_Q0_0_INTRO_96_reg_model LDPC_DEC_ERR_Q0_0_INTRO_96;
    rand LDPC_DEC_ERR_Q0_0_INTRO_97_reg_model LDPC_DEC_ERR_Q0_0_INTRO_97;
    rand LDPC_DEC_ERR_Q0_0_INTRO_98_reg_model LDPC_DEC_ERR_Q0_0_INTRO_98;
    rand LDPC_DEC_ERR_Q0_0_INTRO_99_reg_model LDPC_DEC_ERR_Q0_0_INTRO_99;
    rand LDPC_DEC_ERR_Q0_0_INTRO_100_reg_model LDPC_DEC_ERR_Q0_0_INTRO_100;
    rand LDPC_DEC_ERR_Q0_0_INTRO_101_reg_model LDPC_DEC_ERR_Q0_0_INTRO_101;
    rand LDPC_DEC_ERR_Q0_0_INTRO_102_reg_model LDPC_DEC_ERR_Q0_0_INTRO_102;
    rand LDPC_DEC_ERR_Q0_0_INTRO_103_reg_model LDPC_DEC_ERR_Q0_0_INTRO_103;
    rand LDPC_DEC_ERR_Q0_0_INTRO_104_reg_model LDPC_DEC_ERR_Q0_0_INTRO_104;
    rand LDPC_DEC_ERR_Q0_0_INTRO_105_reg_model LDPC_DEC_ERR_Q0_0_INTRO_105;
    rand LDPC_DEC_ERR_Q0_0_INTRO_106_reg_model LDPC_DEC_ERR_Q0_0_INTRO_106;
    rand LDPC_DEC_ERR_Q0_0_INTRO_107_reg_model LDPC_DEC_ERR_Q0_0_INTRO_107;
    rand LDPC_DEC_ERR_Q0_0_INTRO_108_reg_model LDPC_DEC_ERR_Q0_0_INTRO_108;
    rand LDPC_DEC_ERR_Q0_0_INTRO_109_reg_model LDPC_DEC_ERR_Q0_0_INTRO_109;
    rand LDPC_DEC_ERR_Q0_0_INTRO_110_reg_model LDPC_DEC_ERR_Q0_0_INTRO_110;
    rand LDPC_DEC_ERR_Q0_0_INTRO_111_reg_model LDPC_DEC_ERR_Q0_0_INTRO_111;
    rand LDPC_DEC_ERR_Q0_0_INTRO_112_reg_model LDPC_DEC_ERR_Q0_0_INTRO_112;
    rand LDPC_DEC_ERR_Q0_0_INTRO_113_reg_model LDPC_DEC_ERR_Q0_0_INTRO_113;
    rand LDPC_DEC_ERR_Q0_0_INTRO_114_reg_model LDPC_DEC_ERR_Q0_0_INTRO_114;
    rand LDPC_DEC_ERR_Q0_0_INTRO_115_reg_model LDPC_DEC_ERR_Q0_0_INTRO_115;
    rand LDPC_DEC_ERR_Q0_0_INTRO_116_reg_model LDPC_DEC_ERR_Q0_0_INTRO_116;
    rand LDPC_DEC_ERR_Q0_0_INTRO_117_reg_model LDPC_DEC_ERR_Q0_0_INTRO_117;
    rand LDPC_DEC_ERR_Q0_0_INTRO_118_reg_model LDPC_DEC_ERR_Q0_0_INTRO_118;
    rand LDPC_DEC_ERR_Q0_0_INTRO_119_reg_model LDPC_DEC_ERR_Q0_0_INTRO_119;
    rand LDPC_DEC_ERR_Q0_0_INTRO_120_reg_model LDPC_DEC_ERR_Q0_0_INTRO_120;
    rand LDPC_DEC_ERR_Q0_0_INTRO_121_reg_model LDPC_DEC_ERR_Q0_0_INTRO_121;
    rand LDPC_DEC_ERR_Q0_0_INTRO_122_reg_model LDPC_DEC_ERR_Q0_0_INTRO_122;
    rand LDPC_DEC_ERR_Q0_0_INTRO_123_reg_model LDPC_DEC_ERR_Q0_0_INTRO_123;
    rand LDPC_DEC_ERR_Q0_0_INTRO_124_reg_model LDPC_DEC_ERR_Q0_0_INTRO_124;
    rand LDPC_DEC_ERR_Q0_0_INTRO_125_reg_model LDPC_DEC_ERR_Q0_0_INTRO_125;
    rand LDPC_DEC_ERR_Q0_0_INTRO_126_reg_model LDPC_DEC_ERR_Q0_0_INTRO_126;
    rand LDPC_DEC_ERR_Q0_0_INTRO_127_reg_model LDPC_DEC_ERR_Q0_0_INTRO_127;
    rand LDPC_DEC_ERR_Q0_0_INTRO_128_reg_model LDPC_DEC_ERR_Q0_0_INTRO_128;
    rand LDPC_DEC_ERR_Q0_0_INTRO_129_reg_model LDPC_DEC_ERR_Q0_0_INTRO_129;
    rand LDPC_DEC_ERR_Q0_0_INTRO_130_reg_model LDPC_DEC_ERR_Q0_0_INTRO_130;
    rand LDPC_DEC_ERR_Q0_0_INTRO_131_reg_model LDPC_DEC_ERR_Q0_0_INTRO_131;
    rand LDPC_DEC_ERR_Q0_0_INTRO_132_reg_model LDPC_DEC_ERR_Q0_0_INTRO_132;
    rand LDPC_DEC_ERR_Q0_0_INTRO_133_reg_model LDPC_DEC_ERR_Q0_0_INTRO_133;
    rand LDPC_DEC_ERR_Q0_0_INTRO_134_reg_model LDPC_DEC_ERR_Q0_0_INTRO_134;
    rand LDPC_DEC_ERR_Q0_0_INTRO_135_reg_model LDPC_DEC_ERR_Q0_0_INTRO_135;
    rand LDPC_DEC_ERR_Q0_0_INTRO_136_reg_model LDPC_DEC_ERR_Q0_0_INTRO_136;
    rand LDPC_DEC_ERR_Q0_0_INTRO_137_reg_model LDPC_DEC_ERR_Q0_0_INTRO_137;
    rand LDPC_DEC_ERR_Q0_0_INTRO_138_reg_model LDPC_DEC_ERR_Q0_0_INTRO_138;
    rand LDPC_DEC_ERR_Q0_0_INTRO_139_reg_model LDPC_DEC_ERR_Q0_0_INTRO_139;
    rand LDPC_DEC_ERR_Q0_0_INTRO_140_reg_model LDPC_DEC_ERR_Q0_0_INTRO_140;
    rand LDPC_DEC_ERR_Q0_0_INTRO_141_reg_model LDPC_DEC_ERR_Q0_0_INTRO_141;
    rand LDPC_DEC_ERR_Q0_0_INTRO_142_reg_model LDPC_DEC_ERR_Q0_0_INTRO_142;
    rand LDPC_DEC_ERR_Q0_0_INTRO_143_reg_model LDPC_DEC_ERR_Q0_0_INTRO_143;
    rand LDPC_DEC_ERR_Q0_0_INTRO_144_reg_model LDPC_DEC_ERR_Q0_0_INTRO_144;
    rand LDPC_DEC_ERR_Q0_0_INTRO_145_reg_model LDPC_DEC_ERR_Q0_0_INTRO_145;
    rand LDPC_DEC_ERR_Q0_0_INTRO_146_reg_model LDPC_DEC_ERR_Q0_0_INTRO_146;
    rand LDPC_DEC_ERR_Q0_0_INTRO_147_reg_model LDPC_DEC_ERR_Q0_0_INTRO_147;
    rand LDPC_DEC_ERR_Q0_0_INTRO_148_reg_model LDPC_DEC_ERR_Q0_0_INTRO_148;
    rand LDPC_DEC_ERR_Q0_0_INTRO_149_reg_model LDPC_DEC_ERR_Q0_0_INTRO_149;
    rand LDPC_DEC_ERR_Q0_0_INTRO_150_reg_model LDPC_DEC_ERR_Q0_0_INTRO_150;
    rand LDPC_DEC_ERR_Q0_0_INTRO_151_reg_model LDPC_DEC_ERR_Q0_0_INTRO_151;
    rand LDPC_DEC_ERR_Q0_0_INTRO_152_reg_model LDPC_DEC_ERR_Q0_0_INTRO_152;
    rand LDPC_DEC_ERR_Q0_0_INTRO_153_reg_model LDPC_DEC_ERR_Q0_0_INTRO_153;
    rand LDPC_DEC_ERR_Q0_0_INTRO_154_reg_model LDPC_DEC_ERR_Q0_0_INTRO_154;
    rand LDPC_DEC_ERR_Q0_0_INTRO_155_reg_model LDPC_DEC_ERR_Q0_0_INTRO_155;
    rand LDPC_DEC_ERR_Q0_0_INTRO_156_reg_model LDPC_DEC_ERR_Q0_0_INTRO_156;
    rand LDPC_DEC_ERR_Q0_0_INTRO_157_reg_model LDPC_DEC_ERR_Q0_0_INTRO_157;
    rand LDPC_DEC_ERR_Q0_0_INTRO_158_reg_model LDPC_DEC_ERR_Q0_0_INTRO_158;
    rand LDPC_DEC_ERR_Q0_0_INTRO_159_reg_model LDPC_DEC_ERR_Q0_0_INTRO_159;
    rand LDPC_DEC_ERR_Q0_0_INTRO_160_reg_model LDPC_DEC_ERR_Q0_0_INTRO_160;
    rand LDPC_DEC_ERR_Q0_0_INTRO_161_reg_model LDPC_DEC_ERR_Q0_0_INTRO_161;
    rand LDPC_DEC_ERR_Q0_0_INTRO_162_reg_model LDPC_DEC_ERR_Q0_0_INTRO_162;
    rand LDPC_DEC_ERR_Q0_0_INTRO_163_reg_model LDPC_DEC_ERR_Q0_0_INTRO_163;
    rand LDPC_DEC_ERR_Q0_0_INTRO_164_reg_model LDPC_DEC_ERR_Q0_0_INTRO_164;
    rand LDPC_DEC_ERR_Q0_0_INTRO_165_reg_model LDPC_DEC_ERR_Q0_0_INTRO_165;
    rand LDPC_DEC_ERR_Q0_0_INTRO_166_reg_model LDPC_DEC_ERR_Q0_0_INTRO_166;
    rand LDPC_DEC_ERR_Q0_0_INTRO_167_reg_model LDPC_DEC_ERR_Q0_0_INTRO_167;
    rand LDPC_DEC_ERR_Q0_0_INTRO_168_reg_model LDPC_DEC_ERR_Q0_0_INTRO_168;
    rand LDPC_DEC_ERR_Q0_0_INTRO_169_reg_model LDPC_DEC_ERR_Q0_0_INTRO_169;
    rand LDPC_DEC_ERR_Q0_0_INTRO_170_reg_model LDPC_DEC_ERR_Q0_0_INTRO_170;
    rand LDPC_DEC_ERR_Q0_0_INTRO_171_reg_model LDPC_DEC_ERR_Q0_0_INTRO_171;
    rand LDPC_DEC_ERR_Q0_0_INTRO_172_reg_model LDPC_DEC_ERR_Q0_0_INTRO_172;
    rand LDPC_DEC_ERR_Q0_0_INTRO_173_reg_model LDPC_DEC_ERR_Q0_0_INTRO_173;
    rand LDPC_DEC_ERR_Q0_0_INTRO_174_reg_model LDPC_DEC_ERR_Q0_0_INTRO_174;
    rand LDPC_DEC_ERR_Q0_0_INTRO_175_reg_model LDPC_DEC_ERR_Q0_0_INTRO_175;
    rand LDPC_DEC_ERR_Q0_0_INTRO_176_reg_model LDPC_DEC_ERR_Q0_0_INTRO_176;
    rand LDPC_DEC_ERR_Q0_0_INTRO_177_reg_model LDPC_DEC_ERR_Q0_0_INTRO_177;
    rand LDPC_DEC_ERR_Q0_0_INTRO_178_reg_model LDPC_DEC_ERR_Q0_0_INTRO_178;
    rand LDPC_DEC_ERR_Q0_0_INTRO_179_reg_model LDPC_DEC_ERR_Q0_0_INTRO_179;
    rand LDPC_DEC_ERR_Q0_0_INTRO_180_reg_model LDPC_DEC_ERR_Q0_0_INTRO_180;
    rand LDPC_DEC_ERR_Q0_0_INTRO_181_reg_model LDPC_DEC_ERR_Q0_0_INTRO_181;
    rand LDPC_DEC_ERR_Q0_0_INTRO_182_reg_model LDPC_DEC_ERR_Q0_0_INTRO_182;
    rand LDPC_DEC_ERR_Q0_0_INTRO_183_reg_model LDPC_DEC_ERR_Q0_0_INTRO_183;
    rand LDPC_DEC_ERR_Q0_0_INTRO_184_reg_model LDPC_DEC_ERR_Q0_0_INTRO_184;
    rand LDPC_DEC_ERR_Q0_0_INTRO_185_reg_model LDPC_DEC_ERR_Q0_0_INTRO_185;
    rand LDPC_DEC_ERR_Q0_0_INTRO_186_reg_model LDPC_DEC_ERR_Q0_0_INTRO_186;
    rand LDPC_DEC_ERR_Q0_0_INTRO_187_reg_model LDPC_DEC_ERR_Q0_0_INTRO_187;
    rand LDPC_DEC_ERR_Q0_0_INTRO_188_reg_model LDPC_DEC_ERR_Q0_0_INTRO_188;
    rand LDPC_DEC_ERR_Q0_0_INTRO_189_reg_model LDPC_DEC_ERR_Q0_0_INTRO_189;
    rand LDPC_DEC_ERR_Q0_0_INTRO_190_reg_model LDPC_DEC_ERR_Q0_0_INTRO_190;
    rand LDPC_DEC_ERR_Q0_0_INTRO_191_reg_model LDPC_DEC_ERR_Q0_0_INTRO_191;
    rand LDPC_DEC_ERR_Q0_0_INTRO_192_reg_model LDPC_DEC_ERR_Q0_0_INTRO_192;
    rand LDPC_DEC_ERR_Q0_0_INTRO_193_reg_model LDPC_DEC_ERR_Q0_0_INTRO_193;
    rand LDPC_DEC_ERR_Q0_0_INTRO_194_reg_model LDPC_DEC_ERR_Q0_0_INTRO_194;
    rand LDPC_DEC_ERR_Q0_0_INTRO_195_reg_model LDPC_DEC_ERR_Q0_0_INTRO_195;
    rand LDPC_DEC_ERR_Q0_0_INTRO_196_reg_model LDPC_DEC_ERR_Q0_0_INTRO_196;
    rand LDPC_DEC_ERR_Q0_0_INTRO_197_reg_model LDPC_DEC_ERR_Q0_0_INTRO_197;
    rand LDPC_DEC_ERR_Q0_0_INTRO_198_reg_model LDPC_DEC_ERR_Q0_0_INTRO_198;
    rand LDPC_DEC_ERR_Q0_0_INTRO_199_reg_model LDPC_DEC_ERR_Q0_0_INTRO_199;
    rand LDPC_DEC_ERR_Q0_0_INTRO_200_reg_model LDPC_DEC_ERR_Q0_0_INTRO_200;
    rand LDPC_DEC_ERR_Q0_0_INTRO_201_reg_model LDPC_DEC_ERR_Q0_0_INTRO_201;
    rand LDPC_DEC_ERR_Q0_0_INTRO_202_reg_model LDPC_DEC_ERR_Q0_0_INTRO_202;
    rand LDPC_DEC_ERR_Q0_0_INTRO_203_reg_model LDPC_DEC_ERR_Q0_0_INTRO_203;
    rand LDPC_DEC_ERR_Q0_0_INTRO_204_reg_model LDPC_DEC_ERR_Q0_0_INTRO_204;
    rand LDPC_DEC_ERR_Q0_0_INTRO_205_reg_model LDPC_DEC_ERR_Q0_0_INTRO_205;
    rand LDPC_DEC_ERR_Q0_0_INTRO_206_reg_model LDPC_DEC_ERR_Q0_0_INTRO_206;
    rand LDPC_DEC_ERR_Q0_0_INTRO_207_reg_model LDPC_DEC_ERR_Q0_0_INTRO_207;
    rand LDPC_DEC_ERR_Q0_1_INTRO_0_reg_model LDPC_DEC_ERR_Q0_1_INTRO_0;
    rand LDPC_DEC_ERR_Q0_1_INTRO_1_reg_model LDPC_DEC_ERR_Q0_1_INTRO_1;
    rand LDPC_DEC_ERR_Q0_1_INTRO_2_reg_model LDPC_DEC_ERR_Q0_1_INTRO_2;
    rand LDPC_DEC_ERR_Q0_1_INTRO_3_reg_model LDPC_DEC_ERR_Q0_1_INTRO_3;
    rand LDPC_DEC_ERR_Q0_1_INTRO_4_reg_model LDPC_DEC_ERR_Q0_1_INTRO_4;
    rand LDPC_DEC_ERR_Q0_1_INTRO_5_reg_model LDPC_DEC_ERR_Q0_1_INTRO_5;
    rand LDPC_DEC_ERR_Q0_1_INTRO_6_reg_model LDPC_DEC_ERR_Q0_1_INTRO_6;
    rand LDPC_DEC_ERR_Q0_1_INTRO_7_reg_model LDPC_DEC_ERR_Q0_1_INTRO_7;
    rand LDPC_DEC_ERR_Q0_1_INTRO_8_reg_model LDPC_DEC_ERR_Q0_1_INTRO_8;
    rand LDPC_DEC_ERR_Q0_1_INTRO_9_reg_model LDPC_DEC_ERR_Q0_1_INTRO_9;
    rand LDPC_DEC_ERR_Q0_1_INTRO_10_reg_model LDPC_DEC_ERR_Q0_1_INTRO_10;
    rand LDPC_DEC_ERR_Q0_1_INTRO_11_reg_model LDPC_DEC_ERR_Q0_1_INTRO_11;
    rand LDPC_DEC_ERR_Q0_1_INTRO_12_reg_model LDPC_DEC_ERR_Q0_1_INTRO_12;
    rand LDPC_DEC_ERR_Q0_1_INTRO_13_reg_model LDPC_DEC_ERR_Q0_1_INTRO_13;
    rand LDPC_DEC_ERR_Q0_1_INTRO_14_reg_model LDPC_DEC_ERR_Q0_1_INTRO_14;
    rand LDPC_DEC_ERR_Q0_1_INTRO_15_reg_model LDPC_DEC_ERR_Q0_1_INTRO_15;
    rand LDPC_DEC_ERR_Q0_1_INTRO_16_reg_model LDPC_DEC_ERR_Q0_1_INTRO_16;
    rand LDPC_DEC_ERR_Q0_1_INTRO_17_reg_model LDPC_DEC_ERR_Q0_1_INTRO_17;
    rand LDPC_DEC_ERR_Q0_1_INTRO_18_reg_model LDPC_DEC_ERR_Q0_1_INTRO_18;
    rand LDPC_DEC_ERR_Q0_1_INTRO_19_reg_model LDPC_DEC_ERR_Q0_1_INTRO_19;
    rand LDPC_DEC_ERR_Q0_1_INTRO_20_reg_model LDPC_DEC_ERR_Q0_1_INTRO_20;
    rand LDPC_DEC_ERR_Q0_1_INTRO_21_reg_model LDPC_DEC_ERR_Q0_1_INTRO_21;
    rand LDPC_DEC_ERR_Q0_1_INTRO_22_reg_model LDPC_DEC_ERR_Q0_1_INTRO_22;
    rand LDPC_DEC_ERR_Q0_1_INTRO_23_reg_model LDPC_DEC_ERR_Q0_1_INTRO_23;
    rand LDPC_DEC_ERR_Q0_1_INTRO_24_reg_model LDPC_DEC_ERR_Q0_1_INTRO_24;
    rand LDPC_DEC_ERR_Q0_1_INTRO_25_reg_model LDPC_DEC_ERR_Q0_1_INTRO_25;
    rand LDPC_DEC_ERR_Q0_1_INTRO_26_reg_model LDPC_DEC_ERR_Q0_1_INTRO_26;
    rand LDPC_DEC_ERR_Q0_1_INTRO_27_reg_model LDPC_DEC_ERR_Q0_1_INTRO_27;
    rand LDPC_DEC_ERR_Q0_1_INTRO_28_reg_model LDPC_DEC_ERR_Q0_1_INTRO_28;
    rand LDPC_DEC_ERR_Q0_1_INTRO_29_reg_model LDPC_DEC_ERR_Q0_1_INTRO_29;
    rand LDPC_DEC_ERR_Q0_1_INTRO_30_reg_model LDPC_DEC_ERR_Q0_1_INTRO_30;
    rand LDPC_DEC_ERR_Q0_1_INTRO_31_reg_model LDPC_DEC_ERR_Q0_1_INTRO_31;
    rand LDPC_DEC_ERR_Q0_1_INTRO_32_reg_model LDPC_DEC_ERR_Q0_1_INTRO_32;
    rand LDPC_DEC_ERR_Q0_1_INTRO_33_reg_model LDPC_DEC_ERR_Q0_1_INTRO_33;
    rand LDPC_DEC_ERR_Q0_1_INTRO_34_reg_model LDPC_DEC_ERR_Q0_1_INTRO_34;
    rand LDPC_DEC_ERR_Q0_1_INTRO_35_reg_model LDPC_DEC_ERR_Q0_1_INTRO_35;
    rand LDPC_DEC_ERR_Q0_1_INTRO_36_reg_model LDPC_DEC_ERR_Q0_1_INTRO_36;
    rand LDPC_DEC_ERR_Q0_1_INTRO_37_reg_model LDPC_DEC_ERR_Q0_1_INTRO_37;
    rand LDPC_DEC_ERR_Q0_1_INTRO_38_reg_model LDPC_DEC_ERR_Q0_1_INTRO_38;
    rand LDPC_DEC_ERR_Q0_1_INTRO_39_reg_model LDPC_DEC_ERR_Q0_1_INTRO_39;
    rand LDPC_DEC_ERR_Q0_1_INTRO_40_reg_model LDPC_DEC_ERR_Q0_1_INTRO_40;
    rand LDPC_DEC_ERR_Q0_1_INTRO_41_reg_model LDPC_DEC_ERR_Q0_1_INTRO_41;
    rand LDPC_DEC_ERR_Q0_1_INTRO_42_reg_model LDPC_DEC_ERR_Q0_1_INTRO_42;
    rand LDPC_DEC_ERR_Q0_1_INTRO_43_reg_model LDPC_DEC_ERR_Q0_1_INTRO_43;
    rand LDPC_DEC_ERR_Q0_1_INTRO_44_reg_model LDPC_DEC_ERR_Q0_1_INTRO_44;
    rand LDPC_DEC_ERR_Q0_1_INTRO_45_reg_model LDPC_DEC_ERR_Q0_1_INTRO_45;
    rand LDPC_DEC_ERR_Q0_1_INTRO_46_reg_model LDPC_DEC_ERR_Q0_1_INTRO_46;
    rand LDPC_DEC_ERR_Q0_1_INTRO_47_reg_model LDPC_DEC_ERR_Q0_1_INTRO_47;
    rand LDPC_DEC_ERR_Q0_1_INTRO_48_reg_model LDPC_DEC_ERR_Q0_1_INTRO_48;
    rand LDPC_DEC_ERR_Q0_1_INTRO_49_reg_model LDPC_DEC_ERR_Q0_1_INTRO_49;
    rand LDPC_DEC_ERR_Q0_1_INTRO_50_reg_model LDPC_DEC_ERR_Q0_1_INTRO_50;
    rand LDPC_DEC_ERR_Q0_1_INTRO_51_reg_model LDPC_DEC_ERR_Q0_1_INTRO_51;
    rand LDPC_DEC_ERR_Q0_1_INTRO_52_reg_model LDPC_DEC_ERR_Q0_1_INTRO_52;
    rand LDPC_DEC_ERR_Q0_1_INTRO_53_reg_model LDPC_DEC_ERR_Q0_1_INTRO_53;
    rand LDPC_DEC_ERR_Q0_1_INTRO_54_reg_model LDPC_DEC_ERR_Q0_1_INTRO_54;
    rand LDPC_DEC_ERR_Q0_1_INTRO_55_reg_model LDPC_DEC_ERR_Q0_1_INTRO_55;
    rand LDPC_DEC_ERR_Q0_1_INTRO_56_reg_model LDPC_DEC_ERR_Q0_1_INTRO_56;
    rand LDPC_DEC_ERR_Q0_1_INTRO_57_reg_model LDPC_DEC_ERR_Q0_1_INTRO_57;
    rand LDPC_DEC_ERR_Q0_1_INTRO_58_reg_model LDPC_DEC_ERR_Q0_1_INTRO_58;
    rand LDPC_DEC_ERR_Q0_1_INTRO_59_reg_model LDPC_DEC_ERR_Q0_1_INTRO_59;
    rand LDPC_DEC_ERR_Q0_1_INTRO_60_reg_model LDPC_DEC_ERR_Q0_1_INTRO_60;
    rand LDPC_DEC_ERR_Q0_1_INTRO_61_reg_model LDPC_DEC_ERR_Q0_1_INTRO_61;
    rand LDPC_DEC_ERR_Q0_1_INTRO_62_reg_model LDPC_DEC_ERR_Q0_1_INTRO_62;
    rand LDPC_DEC_ERR_Q0_1_INTRO_63_reg_model LDPC_DEC_ERR_Q0_1_INTRO_63;
    rand LDPC_DEC_ERR_Q0_1_INTRO_64_reg_model LDPC_DEC_ERR_Q0_1_INTRO_64;
    rand LDPC_DEC_ERR_Q0_1_INTRO_65_reg_model LDPC_DEC_ERR_Q0_1_INTRO_65;
    rand LDPC_DEC_ERR_Q0_1_INTRO_66_reg_model LDPC_DEC_ERR_Q0_1_INTRO_66;
    rand LDPC_DEC_ERR_Q0_1_INTRO_67_reg_model LDPC_DEC_ERR_Q0_1_INTRO_67;
    rand LDPC_DEC_ERR_Q0_1_INTRO_68_reg_model LDPC_DEC_ERR_Q0_1_INTRO_68;
    rand LDPC_DEC_ERR_Q0_1_INTRO_69_reg_model LDPC_DEC_ERR_Q0_1_INTRO_69;
    rand LDPC_DEC_ERR_Q0_1_INTRO_70_reg_model LDPC_DEC_ERR_Q0_1_INTRO_70;
    rand LDPC_DEC_ERR_Q0_1_INTRO_71_reg_model LDPC_DEC_ERR_Q0_1_INTRO_71;
    rand LDPC_DEC_ERR_Q0_1_INTRO_72_reg_model LDPC_DEC_ERR_Q0_1_INTRO_72;
    rand LDPC_DEC_ERR_Q0_1_INTRO_73_reg_model LDPC_DEC_ERR_Q0_1_INTRO_73;
    rand LDPC_DEC_ERR_Q0_1_INTRO_74_reg_model LDPC_DEC_ERR_Q0_1_INTRO_74;
    rand LDPC_DEC_ERR_Q0_1_INTRO_75_reg_model LDPC_DEC_ERR_Q0_1_INTRO_75;
    rand LDPC_DEC_ERR_Q0_1_INTRO_76_reg_model LDPC_DEC_ERR_Q0_1_INTRO_76;
    rand LDPC_DEC_ERR_Q0_1_INTRO_77_reg_model LDPC_DEC_ERR_Q0_1_INTRO_77;
    rand LDPC_DEC_ERR_Q0_1_INTRO_78_reg_model LDPC_DEC_ERR_Q0_1_INTRO_78;
    rand LDPC_DEC_ERR_Q0_1_INTRO_79_reg_model LDPC_DEC_ERR_Q0_1_INTRO_79;
    rand LDPC_DEC_ERR_Q0_1_INTRO_80_reg_model LDPC_DEC_ERR_Q0_1_INTRO_80;
    rand LDPC_DEC_ERR_Q0_1_INTRO_81_reg_model LDPC_DEC_ERR_Q0_1_INTRO_81;
    rand LDPC_DEC_ERR_Q0_1_INTRO_82_reg_model LDPC_DEC_ERR_Q0_1_INTRO_82;
    rand LDPC_DEC_ERR_Q0_1_INTRO_83_reg_model LDPC_DEC_ERR_Q0_1_INTRO_83;
    rand LDPC_DEC_ERR_Q0_1_INTRO_84_reg_model LDPC_DEC_ERR_Q0_1_INTRO_84;
    rand LDPC_DEC_ERR_Q0_1_INTRO_85_reg_model LDPC_DEC_ERR_Q0_1_INTRO_85;
    rand LDPC_DEC_ERR_Q0_1_INTRO_86_reg_model LDPC_DEC_ERR_Q0_1_INTRO_86;
    rand LDPC_DEC_ERR_Q0_1_INTRO_87_reg_model LDPC_DEC_ERR_Q0_1_INTRO_87;
    rand LDPC_DEC_ERR_Q0_1_INTRO_88_reg_model LDPC_DEC_ERR_Q0_1_INTRO_88;
    rand LDPC_DEC_ERR_Q0_1_INTRO_89_reg_model LDPC_DEC_ERR_Q0_1_INTRO_89;
    rand LDPC_DEC_ERR_Q0_1_INTRO_90_reg_model LDPC_DEC_ERR_Q0_1_INTRO_90;
    rand LDPC_DEC_ERR_Q0_1_INTRO_91_reg_model LDPC_DEC_ERR_Q0_1_INTRO_91;
    rand LDPC_DEC_ERR_Q0_1_INTRO_92_reg_model LDPC_DEC_ERR_Q0_1_INTRO_92;
    rand LDPC_DEC_ERR_Q0_1_INTRO_93_reg_model LDPC_DEC_ERR_Q0_1_INTRO_93;
    rand LDPC_DEC_ERR_Q0_1_INTRO_94_reg_model LDPC_DEC_ERR_Q0_1_INTRO_94;
    rand LDPC_DEC_ERR_Q0_1_INTRO_95_reg_model LDPC_DEC_ERR_Q0_1_INTRO_95;
    rand LDPC_DEC_ERR_Q0_1_INTRO_96_reg_model LDPC_DEC_ERR_Q0_1_INTRO_96;
    rand LDPC_DEC_ERR_Q0_1_INTRO_97_reg_model LDPC_DEC_ERR_Q0_1_INTRO_97;
    rand LDPC_DEC_ERR_Q0_1_INTRO_98_reg_model LDPC_DEC_ERR_Q0_1_INTRO_98;
    rand LDPC_DEC_ERR_Q0_1_INTRO_99_reg_model LDPC_DEC_ERR_Q0_1_INTRO_99;
    rand LDPC_DEC_ERR_Q0_1_INTRO_100_reg_model LDPC_DEC_ERR_Q0_1_INTRO_100;
    rand LDPC_DEC_ERR_Q0_1_INTRO_101_reg_model LDPC_DEC_ERR_Q0_1_INTRO_101;
    rand LDPC_DEC_ERR_Q0_1_INTRO_102_reg_model LDPC_DEC_ERR_Q0_1_INTRO_102;
    rand LDPC_DEC_ERR_Q0_1_INTRO_103_reg_model LDPC_DEC_ERR_Q0_1_INTRO_103;
    rand LDPC_DEC_ERR_Q0_1_INTRO_104_reg_model LDPC_DEC_ERR_Q0_1_INTRO_104;
    rand LDPC_DEC_ERR_Q0_1_INTRO_105_reg_model LDPC_DEC_ERR_Q0_1_INTRO_105;
    rand LDPC_DEC_ERR_Q0_1_INTRO_106_reg_model LDPC_DEC_ERR_Q0_1_INTRO_106;
    rand LDPC_DEC_ERR_Q0_1_INTRO_107_reg_model LDPC_DEC_ERR_Q0_1_INTRO_107;
    rand LDPC_DEC_ERR_Q0_1_INTRO_108_reg_model LDPC_DEC_ERR_Q0_1_INTRO_108;
    rand LDPC_DEC_ERR_Q0_1_INTRO_109_reg_model LDPC_DEC_ERR_Q0_1_INTRO_109;
    rand LDPC_DEC_ERR_Q0_1_INTRO_110_reg_model LDPC_DEC_ERR_Q0_1_INTRO_110;
    rand LDPC_DEC_ERR_Q0_1_INTRO_111_reg_model LDPC_DEC_ERR_Q0_1_INTRO_111;
    rand LDPC_DEC_ERR_Q0_1_INTRO_112_reg_model LDPC_DEC_ERR_Q0_1_INTRO_112;
    rand LDPC_DEC_ERR_Q0_1_INTRO_113_reg_model LDPC_DEC_ERR_Q0_1_INTRO_113;
    rand LDPC_DEC_ERR_Q0_1_INTRO_114_reg_model LDPC_DEC_ERR_Q0_1_INTRO_114;
    rand LDPC_DEC_ERR_Q0_1_INTRO_115_reg_model LDPC_DEC_ERR_Q0_1_INTRO_115;
    rand LDPC_DEC_ERR_Q0_1_INTRO_116_reg_model LDPC_DEC_ERR_Q0_1_INTRO_116;
    rand LDPC_DEC_ERR_Q0_1_INTRO_117_reg_model LDPC_DEC_ERR_Q0_1_INTRO_117;
    rand LDPC_DEC_ERR_Q0_1_INTRO_118_reg_model LDPC_DEC_ERR_Q0_1_INTRO_118;
    rand LDPC_DEC_ERR_Q0_1_INTRO_119_reg_model LDPC_DEC_ERR_Q0_1_INTRO_119;
    rand LDPC_DEC_ERR_Q0_1_INTRO_120_reg_model LDPC_DEC_ERR_Q0_1_INTRO_120;
    rand LDPC_DEC_ERR_Q0_1_INTRO_121_reg_model LDPC_DEC_ERR_Q0_1_INTRO_121;
    rand LDPC_DEC_ERR_Q0_1_INTRO_122_reg_model LDPC_DEC_ERR_Q0_1_INTRO_122;
    rand LDPC_DEC_ERR_Q0_1_INTRO_123_reg_model LDPC_DEC_ERR_Q0_1_INTRO_123;
    rand LDPC_DEC_ERR_Q0_1_INTRO_124_reg_model LDPC_DEC_ERR_Q0_1_INTRO_124;
    rand LDPC_DEC_ERR_Q0_1_INTRO_125_reg_model LDPC_DEC_ERR_Q0_1_INTRO_125;
    rand LDPC_DEC_ERR_Q0_1_INTRO_126_reg_model LDPC_DEC_ERR_Q0_1_INTRO_126;
    rand LDPC_DEC_ERR_Q0_1_INTRO_127_reg_model LDPC_DEC_ERR_Q0_1_INTRO_127;
    rand LDPC_DEC_ERR_Q0_1_INTRO_128_reg_model LDPC_DEC_ERR_Q0_1_INTRO_128;
    rand LDPC_DEC_ERR_Q0_1_INTRO_129_reg_model LDPC_DEC_ERR_Q0_1_INTRO_129;
    rand LDPC_DEC_ERR_Q0_1_INTRO_130_reg_model LDPC_DEC_ERR_Q0_1_INTRO_130;
    rand LDPC_DEC_ERR_Q0_1_INTRO_131_reg_model LDPC_DEC_ERR_Q0_1_INTRO_131;
    rand LDPC_DEC_ERR_Q0_1_INTRO_132_reg_model LDPC_DEC_ERR_Q0_1_INTRO_132;
    rand LDPC_DEC_ERR_Q0_1_INTRO_133_reg_model LDPC_DEC_ERR_Q0_1_INTRO_133;
    rand LDPC_DEC_ERR_Q0_1_INTRO_134_reg_model LDPC_DEC_ERR_Q0_1_INTRO_134;
    rand LDPC_DEC_ERR_Q0_1_INTRO_135_reg_model LDPC_DEC_ERR_Q0_1_INTRO_135;
    rand LDPC_DEC_ERR_Q0_1_INTRO_136_reg_model LDPC_DEC_ERR_Q0_1_INTRO_136;
    rand LDPC_DEC_ERR_Q0_1_INTRO_137_reg_model LDPC_DEC_ERR_Q0_1_INTRO_137;
    rand LDPC_DEC_ERR_Q0_1_INTRO_138_reg_model LDPC_DEC_ERR_Q0_1_INTRO_138;
    rand LDPC_DEC_ERR_Q0_1_INTRO_139_reg_model LDPC_DEC_ERR_Q0_1_INTRO_139;
    rand LDPC_DEC_ERR_Q0_1_INTRO_140_reg_model LDPC_DEC_ERR_Q0_1_INTRO_140;
    rand LDPC_DEC_ERR_Q0_1_INTRO_141_reg_model LDPC_DEC_ERR_Q0_1_INTRO_141;
    rand LDPC_DEC_ERR_Q0_1_INTRO_142_reg_model LDPC_DEC_ERR_Q0_1_INTRO_142;
    rand LDPC_DEC_ERR_Q0_1_INTRO_143_reg_model LDPC_DEC_ERR_Q0_1_INTRO_143;
    rand LDPC_DEC_ERR_Q0_1_INTRO_144_reg_model LDPC_DEC_ERR_Q0_1_INTRO_144;
    rand LDPC_DEC_ERR_Q0_1_INTRO_145_reg_model LDPC_DEC_ERR_Q0_1_INTRO_145;
    rand LDPC_DEC_ERR_Q0_1_INTRO_146_reg_model LDPC_DEC_ERR_Q0_1_INTRO_146;
    rand LDPC_DEC_ERR_Q0_1_INTRO_147_reg_model LDPC_DEC_ERR_Q0_1_INTRO_147;
    rand LDPC_DEC_ERR_Q0_1_INTRO_148_reg_model LDPC_DEC_ERR_Q0_1_INTRO_148;
    rand LDPC_DEC_ERR_Q0_1_INTRO_149_reg_model LDPC_DEC_ERR_Q0_1_INTRO_149;
    rand LDPC_DEC_ERR_Q0_1_INTRO_150_reg_model LDPC_DEC_ERR_Q0_1_INTRO_150;
    rand LDPC_DEC_ERR_Q0_1_INTRO_151_reg_model LDPC_DEC_ERR_Q0_1_INTRO_151;
    rand LDPC_DEC_ERR_Q0_1_INTRO_152_reg_model LDPC_DEC_ERR_Q0_1_INTRO_152;
    rand LDPC_DEC_ERR_Q0_1_INTRO_153_reg_model LDPC_DEC_ERR_Q0_1_INTRO_153;
    rand LDPC_DEC_ERR_Q0_1_INTRO_154_reg_model LDPC_DEC_ERR_Q0_1_INTRO_154;
    rand LDPC_DEC_ERR_Q0_1_INTRO_155_reg_model LDPC_DEC_ERR_Q0_1_INTRO_155;
    rand LDPC_DEC_ERR_Q0_1_INTRO_156_reg_model LDPC_DEC_ERR_Q0_1_INTRO_156;
    rand LDPC_DEC_ERR_Q0_1_INTRO_157_reg_model LDPC_DEC_ERR_Q0_1_INTRO_157;
    rand LDPC_DEC_ERR_Q0_1_INTRO_158_reg_model LDPC_DEC_ERR_Q0_1_INTRO_158;
    rand LDPC_DEC_ERR_Q0_1_INTRO_159_reg_model LDPC_DEC_ERR_Q0_1_INTRO_159;
    rand LDPC_DEC_ERR_Q0_1_INTRO_160_reg_model LDPC_DEC_ERR_Q0_1_INTRO_160;
    rand LDPC_DEC_ERR_Q0_1_INTRO_161_reg_model LDPC_DEC_ERR_Q0_1_INTRO_161;
    rand LDPC_DEC_ERR_Q0_1_INTRO_162_reg_model LDPC_DEC_ERR_Q0_1_INTRO_162;
    rand LDPC_DEC_ERR_Q0_1_INTRO_163_reg_model LDPC_DEC_ERR_Q0_1_INTRO_163;
    rand LDPC_DEC_ERR_Q0_1_INTRO_164_reg_model LDPC_DEC_ERR_Q0_1_INTRO_164;
    rand LDPC_DEC_ERR_Q0_1_INTRO_165_reg_model LDPC_DEC_ERR_Q0_1_INTRO_165;
    rand LDPC_DEC_ERR_Q0_1_INTRO_166_reg_model LDPC_DEC_ERR_Q0_1_INTRO_166;
    rand LDPC_DEC_ERR_Q0_1_INTRO_167_reg_model LDPC_DEC_ERR_Q0_1_INTRO_167;
    rand LDPC_DEC_ERR_Q0_1_INTRO_168_reg_model LDPC_DEC_ERR_Q0_1_INTRO_168;
    rand LDPC_DEC_ERR_Q0_1_INTRO_169_reg_model LDPC_DEC_ERR_Q0_1_INTRO_169;
    rand LDPC_DEC_ERR_Q0_1_INTRO_170_reg_model LDPC_DEC_ERR_Q0_1_INTRO_170;
    rand LDPC_DEC_ERR_Q0_1_INTRO_171_reg_model LDPC_DEC_ERR_Q0_1_INTRO_171;
    rand LDPC_DEC_ERR_Q0_1_INTRO_172_reg_model LDPC_DEC_ERR_Q0_1_INTRO_172;
    rand LDPC_DEC_ERR_Q0_1_INTRO_173_reg_model LDPC_DEC_ERR_Q0_1_INTRO_173;
    rand LDPC_DEC_ERR_Q0_1_INTRO_174_reg_model LDPC_DEC_ERR_Q0_1_INTRO_174;
    rand LDPC_DEC_ERR_Q0_1_INTRO_175_reg_model LDPC_DEC_ERR_Q0_1_INTRO_175;
    rand LDPC_DEC_ERR_Q0_1_INTRO_176_reg_model LDPC_DEC_ERR_Q0_1_INTRO_176;
    rand LDPC_DEC_ERR_Q0_1_INTRO_177_reg_model LDPC_DEC_ERR_Q0_1_INTRO_177;
    rand LDPC_DEC_ERR_Q0_1_INTRO_178_reg_model LDPC_DEC_ERR_Q0_1_INTRO_178;
    rand LDPC_DEC_ERR_Q0_1_INTRO_179_reg_model LDPC_DEC_ERR_Q0_1_INTRO_179;
    rand LDPC_DEC_ERR_Q0_1_INTRO_180_reg_model LDPC_DEC_ERR_Q0_1_INTRO_180;
    rand LDPC_DEC_ERR_Q0_1_INTRO_181_reg_model LDPC_DEC_ERR_Q0_1_INTRO_181;
    rand LDPC_DEC_ERR_Q0_1_INTRO_182_reg_model LDPC_DEC_ERR_Q0_1_INTRO_182;
    rand LDPC_DEC_ERR_Q0_1_INTRO_183_reg_model LDPC_DEC_ERR_Q0_1_INTRO_183;
    rand LDPC_DEC_ERR_Q0_1_INTRO_184_reg_model LDPC_DEC_ERR_Q0_1_INTRO_184;
    rand LDPC_DEC_ERR_Q0_1_INTRO_185_reg_model LDPC_DEC_ERR_Q0_1_INTRO_185;
    rand LDPC_DEC_ERR_Q0_1_INTRO_186_reg_model LDPC_DEC_ERR_Q0_1_INTRO_186;
    rand LDPC_DEC_ERR_Q0_1_INTRO_187_reg_model LDPC_DEC_ERR_Q0_1_INTRO_187;
    rand LDPC_DEC_ERR_Q0_1_INTRO_188_reg_model LDPC_DEC_ERR_Q0_1_INTRO_188;
    rand LDPC_DEC_ERR_Q0_1_INTRO_189_reg_model LDPC_DEC_ERR_Q0_1_INTRO_189;
    rand LDPC_DEC_ERR_Q0_1_INTRO_190_reg_model LDPC_DEC_ERR_Q0_1_INTRO_190;
    rand LDPC_DEC_ERR_Q0_1_INTRO_191_reg_model LDPC_DEC_ERR_Q0_1_INTRO_191;
    rand LDPC_DEC_ERR_Q0_1_INTRO_192_reg_model LDPC_DEC_ERR_Q0_1_INTRO_192;
    rand LDPC_DEC_ERR_Q0_1_INTRO_193_reg_model LDPC_DEC_ERR_Q0_1_INTRO_193;
    rand LDPC_DEC_ERR_Q0_1_INTRO_194_reg_model LDPC_DEC_ERR_Q0_1_INTRO_194;
    rand LDPC_DEC_ERR_Q0_1_INTRO_195_reg_model LDPC_DEC_ERR_Q0_1_INTRO_195;
    rand LDPC_DEC_ERR_Q0_1_INTRO_196_reg_model LDPC_DEC_ERR_Q0_1_INTRO_196;
    rand LDPC_DEC_ERR_Q0_1_INTRO_197_reg_model LDPC_DEC_ERR_Q0_1_INTRO_197;
    rand LDPC_DEC_ERR_Q0_1_INTRO_198_reg_model LDPC_DEC_ERR_Q0_1_INTRO_198;
    rand LDPC_DEC_ERR_Q0_1_INTRO_199_reg_model LDPC_DEC_ERR_Q0_1_INTRO_199;
    rand LDPC_DEC_ERR_Q0_1_INTRO_200_reg_model LDPC_DEC_ERR_Q0_1_INTRO_200;
    rand LDPC_DEC_ERR_Q0_1_INTRO_201_reg_model LDPC_DEC_ERR_Q0_1_INTRO_201;
    rand LDPC_DEC_ERR_Q0_1_INTRO_202_reg_model LDPC_DEC_ERR_Q0_1_INTRO_202;
    rand LDPC_DEC_ERR_Q0_1_INTRO_203_reg_model LDPC_DEC_ERR_Q0_1_INTRO_203;
    rand LDPC_DEC_ERR_Q0_1_INTRO_204_reg_model LDPC_DEC_ERR_Q0_1_INTRO_204;
    rand LDPC_DEC_ERR_Q0_1_INTRO_205_reg_model LDPC_DEC_ERR_Q0_1_INTRO_205;
    rand LDPC_DEC_ERR_Q0_1_INTRO_206_reg_model LDPC_DEC_ERR_Q0_1_INTRO_206;
    rand LDPC_DEC_ERR_Q0_1_INTRO_207_reg_model LDPC_DEC_ERR_Q0_1_INTRO_207;
    rand LDPC_DEC_ERR_INTRODUCED_reg_model LDPC_DEC_ERR_INTRODUCED;
    rand LDPC_DEC_CODEWRD_IN_q0_0_0_reg_model LDPC_DEC_CODEWRD_IN_q0_0_0;
    rand LDPC_DEC_CODEWRD_IN_q0_0_1_reg_model LDPC_DEC_CODEWRD_IN_q0_0_1;
    rand LDPC_DEC_CODEWRD_IN_q0_0_2_reg_model LDPC_DEC_CODEWRD_IN_q0_0_2;
    rand LDPC_DEC_CODEWRD_IN_q0_0_3_reg_model LDPC_DEC_CODEWRD_IN_q0_0_3;
    rand LDPC_DEC_CODEWRD_IN_q0_0_4_reg_model LDPC_DEC_CODEWRD_IN_q0_0_4;
    rand LDPC_DEC_CODEWRD_IN_q0_0_5_reg_model LDPC_DEC_CODEWRD_IN_q0_0_5;
    rand LDPC_DEC_CODEWRD_IN_q0_0_6_reg_model LDPC_DEC_CODEWRD_IN_q0_0_6;
    rand LDPC_DEC_CODEWRD_IN_q0_0_7_reg_model LDPC_DEC_CODEWRD_IN_q0_0_7;
    rand LDPC_DEC_CODEWRD_IN_q0_0_8_reg_model LDPC_DEC_CODEWRD_IN_q0_0_8;
    rand LDPC_DEC_CODEWRD_IN_q0_0_9_reg_model LDPC_DEC_CODEWRD_IN_q0_0_9;
    rand LDPC_DEC_CODEWRD_IN_q0_0_10_reg_model LDPC_DEC_CODEWRD_IN_q0_0_10;
    rand LDPC_DEC_CODEWRD_IN_q0_0_11_reg_model LDPC_DEC_CODEWRD_IN_q0_0_11;
    rand LDPC_DEC_CODEWRD_IN_q0_0_12_reg_model LDPC_DEC_CODEWRD_IN_q0_0_12;
    rand LDPC_DEC_CODEWRD_IN_q0_0_13_reg_model LDPC_DEC_CODEWRD_IN_q0_0_13;
    rand LDPC_DEC_CODEWRD_IN_q0_0_14_reg_model LDPC_DEC_CODEWRD_IN_q0_0_14;
    rand LDPC_DEC_CODEWRD_IN_q0_0_15_reg_model LDPC_DEC_CODEWRD_IN_q0_0_15;
    rand LDPC_DEC_CODEWRD_IN_q0_0_16_reg_model LDPC_DEC_CODEWRD_IN_q0_0_16;
    rand LDPC_DEC_CODEWRD_IN_q0_0_17_reg_model LDPC_DEC_CODEWRD_IN_q0_0_17;
    rand LDPC_DEC_CODEWRD_IN_q0_0_18_reg_model LDPC_DEC_CODEWRD_IN_q0_0_18;
    rand LDPC_DEC_CODEWRD_IN_q0_0_19_reg_model LDPC_DEC_CODEWRD_IN_q0_0_19;
    rand LDPC_DEC_CODEWRD_IN_q0_0_20_reg_model LDPC_DEC_CODEWRD_IN_q0_0_20;
    rand LDPC_DEC_CODEWRD_IN_q0_0_21_reg_model LDPC_DEC_CODEWRD_IN_q0_0_21;
    rand LDPC_DEC_CODEWRD_IN_q0_0_22_reg_model LDPC_DEC_CODEWRD_IN_q0_0_22;
    rand LDPC_DEC_CODEWRD_IN_q0_0_23_reg_model LDPC_DEC_CODEWRD_IN_q0_0_23;
    rand LDPC_DEC_CODEWRD_IN_q0_0_24_reg_model LDPC_DEC_CODEWRD_IN_q0_0_24;
    rand LDPC_DEC_CODEWRD_IN_q0_0_25_reg_model LDPC_DEC_CODEWRD_IN_q0_0_25;
    rand LDPC_DEC_CODEWRD_IN_q0_0_26_reg_model LDPC_DEC_CODEWRD_IN_q0_0_26;
    rand LDPC_DEC_CODEWRD_IN_q0_0_27_reg_model LDPC_DEC_CODEWRD_IN_q0_0_27;
    rand LDPC_DEC_CODEWRD_IN_q0_0_28_reg_model LDPC_DEC_CODEWRD_IN_q0_0_28;
    rand LDPC_DEC_CODEWRD_IN_q0_0_29_reg_model LDPC_DEC_CODEWRD_IN_q0_0_29;
    rand LDPC_DEC_CODEWRD_IN_q0_0_30_reg_model LDPC_DEC_CODEWRD_IN_q0_0_30;
    rand LDPC_DEC_CODEWRD_IN_q0_0_31_reg_model LDPC_DEC_CODEWRD_IN_q0_0_31;
    rand LDPC_DEC_CODEWRD_IN_q0_0_32_reg_model LDPC_DEC_CODEWRD_IN_q0_0_32;
    rand LDPC_DEC_CODEWRD_IN_q0_0_33_reg_model LDPC_DEC_CODEWRD_IN_q0_0_33;
    rand LDPC_DEC_CODEWRD_IN_q0_0_34_reg_model LDPC_DEC_CODEWRD_IN_q0_0_34;
    rand LDPC_DEC_CODEWRD_IN_q0_0_35_reg_model LDPC_DEC_CODEWRD_IN_q0_0_35;
    rand LDPC_DEC_CODEWRD_IN_q0_0_36_reg_model LDPC_DEC_CODEWRD_IN_q0_0_36;
    rand LDPC_DEC_CODEWRD_IN_q0_0_37_reg_model LDPC_DEC_CODEWRD_IN_q0_0_37;
    rand LDPC_DEC_CODEWRD_IN_q0_0_38_reg_model LDPC_DEC_CODEWRD_IN_q0_0_38;
    rand LDPC_DEC_CODEWRD_IN_q0_0_39_reg_model LDPC_DEC_CODEWRD_IN_q0_0_39;
    rand LDPC_DEC_CODEWRD_IN_q0_0_40_reg_model LDPC_DEC_CODEWRD_IN_q0_0_40;
    rand LDPC_DEC_CODEWRD_IN_q0_0_41_reg_model LDPC_DEC_CODEWRD_IN_q0_0_41;
    rand LDPC_DEC_CODEWRD_IN_q0_0_42_reg_model LDPC_DEC_CODEWRD_IN_q0_0_42;
    rand LDPC_DEC_CODEWRD_IN_q0_0_43_reg_model LDPC_DEC_CODEWRD_IN_q0_0_43;
    rand LDPC_DEC_CODEWRD_IN_q0_0_44_reg_model LDPC_DEC_CODEWRD_IN_q0_0_44;
    rand LDPC_DEC_CODEWRD_IN_q0_0_45_reg_model LDPC_DEC_CODEWRD_IN_q0_0_45;
    rand LDPC_DEC_CODEWRD_IN_q0_0_46_reg_model LDPC_DEC_CODEWRD_IN_q0_0_46;
    rand LDPC_DEC_CODEWRD_IN_q0_0_47_reg_model LDPC_DEC_CODEWRD_IN_q0_0_47;
    rand LDPC_DEC_CODEWRD_IN_q0_0_48_reg_model LDPC_DEC_CODEWRD_IN_q0_0_48;
    rand LDPC_DEC_CODEWRD_IN_q0_0_49_reg_model LDPC_DEC_CODEWRD_IN_q0_0_49;
    rand LDPC_DEC_CODEWRD_IN_q0_0_50_reg_model LDPC_DEC_CODEWRD_IN_q0_0_50;
    rand LDPC_DEC_CODEWRD_IN_q0_0_51_reg_model LDPC_DEC_CODEWRD_IN_q0_0_51;
    rand LDPC_DEC_CODEWRD_IN_q0_0_52_reg_model LDPC_DEC_CODEWRD_IN_q0_0_52;
    rand LDPC_DEC_CODEWRD_IN_q0_0_53_reg_model LDPC_DEC_CODEWRD_IN_q0_0_53;
    rand LDPC_DEC_CODEWRD_IN_q0_0_54_reg_model LDPC_DEC_CODEWRD_IN_q0_0_54;
    rand LDPC_DEC_CODEWRD_IN_q0_0_55_reg_model LDPC_DEC_CODEWRD_IN_q0_0_55;
    rand LDPC_DEC_CODEWRD_IN_q0_0_56_reg_model LDPC_DEC_CODEWRD_IN_q0_0_56;
    rand LDPC_DEC_CODEWRD_IN_q0_0_57_reg_model LDPC_DEC_CODEWRD_IN_q0_0_57;
    rand LDPC_DEC_CODEWRD_IN_q0_0_58_reg_model LDPC_DEC_CODEWRD_IN_q0_0_58;
    rand LDPC_DEC_CODEWRD_IN_q0_0_59_reg_model LDPC_DEC_CODEWRD_IN_q0_0_59;
    rand LDPC_DEC_CODEWRD_IN_q0_0_60_reg_model LDPC_DEC_CODEWRD_IN_q0_0_60;
    rand LDPC_DEC_CODEWRD_IN_q0_0_61_reg_model LDPC_DEC_CODEWRD_IN_q0_0_61;
    rand LDPC_DEC_CODEWRD_IN_q0_0_62_reg_model LDPC_DEC_CODEWRD_IN_q0_0_62;
    rand LDPC_DEC_CODEWRD_IN_q0_0_63_reg_model LDPC_DEC_CODEWRD_IN_q0_0_63;
    rand LDPC_DEC_CODEWRD_IN_q0_0_64_reg_model LDPC_DEC_CODEWRD_IN_q0_0_64;
    rand LDPC_DEC_CODEWRD_IN_q0_0_65_reg_model LDPC_DEC_CODEWRD_IN_q0_0_65;
    rand LDPC_DEC_CODEWRD_IN_q0_0_66_reg_model LDPC_DEC_CODEWRD_IN_q0_0_66;
    rand LDPC_DEC_CODEWRD_IN_q0_0_67_reg_model LDPC_DEC_CODEWRD_IN_q0_0_67;
    rand LDPC_DEC_CODEWRD_IN_q0_0_68_reg_model LDPC_DEC_CODEWRD_IN_q0_0_68;
    rand LDPC_DEC_CODEWRD_IN_q0_0_69_reg_model LDPC_DEC_CODEWRD_IN_q0_0_69;
    rand LDPC_DEC_CODEWRD_IN_q0_0_70_reg_model LDPC_DEC_CODEWRD_IN_q0_0_70;
    rand LDPC_DEC_CODEWRD_IN_q0_0_71_reg_model LDPC_DEC_CODEWRD_IN_q0_0_71;
    rand LDPC_DEC_CODEWRD_IN_q0_0_72_reg_model LDPC_DEC_CODEWRD_IN_q0_0_72;
    rand LDPC_DEC_CODEWRD_IN_q0_0_73_reg_model LDPC_DEC_CODEWRD_IN_q0_0_73;
    rand LDPC_DEC_CODEWRD_IN_q0_0_74_reg_model LDPC_DEC_CODEWRD_IN_q0_0_74;
    rand LDPC_DEC_CODEWRD_IN_q0_0_75_reg_model LDPC_DEC_CODEWRD_IN_q0_0_75;
    rand LDPC_DEC_CODEWRD_IN_q0_0_76_reg_model LDPC_DEC_CODEWRD_IN_q0_0_76;
    rand LDPC_DEC_CODEWRD_IN_q0_0_77_reg_model LDPC_DEC_CODEWRD_IN_q0_0_77;
    rand LDPC_DEC_CODEWRD_IN_q0_0_78_reg_model LDPC_DEC_CODEWRD_IN_q0_0_78;
    rand LDPC_DEC_CODEWRD_IN_q0_0_79_reg_model LDPC_DEC_CODEWRD_IN_q0_0_79;
    rand LDPC_DEC_CODEWRD_IN_q0_0_80_reg_model LDPC_DEC_CODEWRD_IN_q0_0_80;
    rand LDPC_DEC_CODEWRD_IN_q0_0_81_reg_model LDPC_DEC_CODEWRD_IN_q0_0_81;
    rand LDPC_DEC_CODEWRD_IN_q0_0_82_reg_model LDPC_DEC_CODEWRD_IN_q0_0_82;
    rand LDPC_DEC_CODEWRD_IN_q0_0_83_reg_model LDPC_DEC_CODEWRD_IN_q0_0_83;
    rand LDPC_DEC_CODEWRD_IN_q0_0_84_reg_model LDPC_DEC_CODEWRD_IN_q0_0_84;
    rand LDPC_DEC_CODEWRD_IN_q0_0_85_reg_model LDPC_DEC_CODEWRD_IN_q0_0_85;
    rand LDPC_DEC_CODEWRD_IN_q0_0_86_reg_model LDPC_DEC_CODEWRD_IN_q0_0_86;
    rand LDPC_DEC_CODEWRD_IN_q0_0_87_reg_model LDPC_DEC_CODEWRD_IN_q0_0_87;
    rand LDPC_DEC_CODEWRD_IN_q0_0_88_reg_model LDPC_DEC_CODEWRD_IN_q0_0_88;
    rand LDPC_DEC_CODEWRD_IN_q0_0_89_reg_model LDPC_DEC_CODEWRD_IN_q0_0_89;
    rand LDPC_DEC_CODEWRD_IN_q0_0_90_reg_model LDPC_DEC_CODEWRD_IN_q0_0_90;
    rand LDPC_DEC_CODEWRD_IN_q0_0_91_reg_model LDPC_DEC_CODEWRD_IN_q0_0_91;
    rand LDPC_DEC_CODEWRD_IN_q0_0_92_reg_model LDPC_DEC_CODEWRD_IN_q0_0_92;
    rand LDPC_DEC_CODEWRD_IN_q0_0_93_reg_model LDPC_DEC_CODEWRD_IN_q0_0_93;
    rand LDPC_DEC_CODEWRD_IN_q0_0_94_reg_model LDPC_DEC_CODEWRD_IN_q0_0_94;
    rand LDPC_DEC_CODEWRD_IN_q0_0_95_reg_model LDPC_DEC_CODEWRD_IN_q0_0_95;
    rand LDPC_DEC_CODEWRD_IN_q0_0_96_reg_model LDPC_DEC_CODEWRD_IN_q0_0_96;
    rand LDPC_DEC_CODEWRD_IN_q0_0_97_reg_model LDPC_DEC_CODEWRD_IN_q0_0_97;
    rand LDPC_DEC_CODEWRD_IN_q0_0_98_reg_model LDPC_DEC_CODEWRD_IN_q0_0_98;
    rand LDPC_DEC_CODEWRD_IN_q0_0_99_reg_model LDPC_DEC_CODEWRD_IN_q0_0_99;
    rand LDPC_DEC_CODEWRD_IN_q0_0_100_reg_model LDPC_DEC_CODEWRD_IN_q0_0_100;
    rand LDPC_DEC_CODEWRD_IN_q0_0_101_reg_model LDPC_DEC_CODEWRD_IN_q0_0_101;
    rand LDPC_DEC_CODEWRD_IN_q0_0_102_reg_model LDPC_DEC_CODEWRD_IN_q0_0_102;
    rand LDPC_DEC_CODEWRD_IN_q0_0_103_reg_model LDPC_DEC_CODEWRD_IN_q0_0_103;
    rand LDPC_DEC_CODEWRD_IN_q0_0_104_reg_model LDPC_DEC_CODEWRD_IN_q0_0_104;
    rand LDPC_DEC_CODEWRD_IN_q0_0_105_reg_model LDPC_DEC_CODEWRD_IN_q0_0_105;
    rand LDPC_DEC_CODEWRD_IN_q0_0_106_reg_model LDPC_DEC_CODEWRD_IN_q0_0_106;
    rand LDPC_DEC_CODEWRD_IN_q0_0_107_reg_model LDPC_DEC_CODEWRD_IN_q0_0_107;
    rand LDPC_DEC_CODEWRD_IN_q0_0_108_reg_model LDPC_DEC_CODEWRD_IN_q0_0_108;
    rand LDPC_DEC_CODEWRD_IN_q0_0_109_reg_model LDPC_DEC_CODEWRD_IN_q0_0_109;
    rand LDPC_DEC_CODEWRD_IN_q0_0_110_reg_model LDPC_DEC_CODEWRD_IN_q0_0_110;
    rand LDPC_DEC_CODEWRD_IN_q0_0_111_reg_model LDPC_DEC_CODEWRD_IN_q0_0_111;
    rand LDPC_DEC_CODEWRD_IN_q0_0_112_reg_model LDPC_DEC_CODEWRD_IN_q0_0_112;
    rand LDPC_DEC_CODEWRD_IN_q0_0_113_reg_model LDPC_DEC_CODEWRD_IN_q0_0_113;
    rand LDPC_DEC_CODEWRD_IN_q0_0_114_reg_model LDPC_DEC_CODEWRD_IN_q0_0_114;
    rand LDPC_DEC_CODEWRD_IN_q0_0_115_reg_model LDPC_DEC_CODEWRD_IN_q0_0_115;
    rand LDPC_DEC_CODEWRD_IN_q0_0_116_reg_model LDPC_DEC_CODEWRD_IN_q0_0_116;
    rand LDPC_DEC_CODEWRD_IN_q0_0_117_reg_model LDPC_DEC_CODEWRD_IN_q0_0_117;
    rand LDPC_DEC_CODEWRD_IN_q0_0_118_reg_model LDPC_DEC_CODEWRD_IN_q0_0_118;
    rand LDPC_DEC_CODEWRD_IN_q0_0_119_reg_model LDPC_DEC_CODEWRD_IN_q0_0_119;
    rand LDPC_DEC_CODEWRD_IN_q0_0_120_reg_model LDPC_DEC_CODEWRD_IN_q0_0_120;
    rand LDPC_DEC_CODEWRD_IN_q0_0_121_reg_model LDPC_DEC_CODEWRD_IN_q0_0_121;
    rand LDPC_DEC_CODEWRD_IN_q0_0_122_reg_model LDPC_DEC_CODEWRD_IN_q0_0_122;
    rand LDPC_DEC_CODEWRD_IN_q0_0_123_reg_model LDPC_DEC_CODEWRD_IN_q0_0_123;
    rand LDPC_DEC_CODEWRD_IN_q0_0_124_reg_model LDPC_DEC_CODEWRD_IN_q0_0_124;
    rand LDPC_DEC_CODEWRD_IN_q0_0_125_reg_model LDPC_DEC_CODEWRD_IN_q0_0_125;
    rand LDPC_DEC_CODEWRD_IN_q0_0_126_reg_model LDPC_DEC_CODEWRD_IN_q0_0_126;
    rand LDPC_DEC_CODEWRD_IN_q0_0_127_reg_model LDPC_DEC_CODEWRD_IN_q0_0_127;
    rand LDPC_DEC_CODEWRD_IN_q0_0_128_reg_model LDPC_DEC_CODEWRD_IN_q0_0_128;
    rand LDPC_DEC_CODEWRD_IN_q0_0_129_reg_model LDPC_DEC_CODEWRD_IN_q0_0_129;
    rand LDPC_DEC_CODEWRD_IN_q0_0_130_reg_model LDPC_DEC_CODEWRD_IN_q0_0_130;
    rand LDPC_DEC_CODEWRD_IN_q0_0_131_reg_model LDPC_DEC_CODEWRD_IN_q0_0_131;
    rand LDPC_DEC_CODEWRD_IN_q0_0_132_reg_model LDPC_DEC_CODEWRD_IN_q0_0_132;
    rand LDPC_DEC_CODEWRD_IN_q0_0_133_reg_model LDPC_DEC_CODEWRD_IN_q0_0_133;
    rand LDPC_DEC_CODEWRD_IN_q0_0_134_reg_model LDPC_DEC_CODEWRD_IN_q0_0_134;
    rand LDPC_DEC_CODEWRD_IN_q0_0_135_reg_model LDPC_DEC_CODEWRD_IN_q0_0_135;
    rand LDPC_DEC_CODEWRD_IN_q0_0_136_reg_model LDPC_DEC_CODEWRD_IN_q0_0_136;
    rand LDPC_DEC_CODEWRD_IN_q0_0_137_reg_model LDPC_DEC_CODEWRD_IN_q0_0_137;
    rand LDPC_DEC_CODEWRD_IN_q0_0_138_reg_model LDPC_DEC_CODEWRD_IN_q0_0_138;
    rand LDPC_DEC_CODEWRD_IN_q0_0_139_reg_model LDPC_DEC_CODEWRD_IN_q0_0_139;
    rand LDPC_DEC_CODEWRD_IN_q0_0_140_reg_model LDPC_DEC_CODEWRD_IN_q0_0_140;
    rand LDPC_DEC_CODEWRD_IN_q0_0_141_reg_model LDPC_DEC_CODEWRD_IN_q0_0_141;
    rand LDPC_DEC_CODEWRD_IN_q0_0_142_reg_model LDPC_DEC_CODEWRD_IN_q0_0_142;
    rand LDPC_DEC_CODEWRD_IN_q0_0_143_reg_model LDPC_DEC_CODEWRD_IN_q0_0_143;
    rand LDPC_DEC_CODEWRD_IN_q0_0_144_reg_model LDPC_DEC_CODEWRD_IN_q0_0_144;
    rand LDPC_DEC_CODEWRD_IN_q0_0_145_reg_model LDPC_DEC_CODEWRD_IN_q0_0_145;
    rand LDPC_DEC_CODEWRD_IN_q0_0_146_reg_model LDPC_DEC_CODEWRD_IN_q0_0_146;
    rand LDPC_DEC_CODEWRD_IN_q0_0_147_reg_model LDPC_DEC_CODEWRD_IN_q0_0_147;
    rand LDPC_DEC_CODEWRD_IN_q0_0_148_reg_model LDPC_DEC_CODEWRD_IN_q0_0_148;
    rand LDPC_DEC_CODEWRD_IN_q0_0_149_reg_model LDPC_DEC_CODEWRD_IN_q0_0_149;
    rand LDPC_DEC_CODEWRD_IN_q0_0_150_reg_model LDPC_DEC_CODEWRD_IN_q0_0_150;
    rand LDPC_DEC_CODEWRD_IN_q0_0_151_reg_model LDPC_DEC_CODEWRD_IN_q0_0_151;
    rand LDPC_DEC_CODEWRD_IN_q0_0_152_reg_model LDPC_DEC_CODEWRD_IN_q0_0_152;
    rand LDPC_DEC_CODEWRD_IN_q0_0_153_reg_model LDPC_DEC_CODEWRD_IN_q0_0_153;
    rand LDPC_DEC_CODEWRD_IN_q0_0_154_reg_model LDPC_DEC_CODEWRD_IN_q0_0_154;
    rand LDPC_DEC_CODEWRD_IN_q0_0_155_reg_model LDPC_DEC_CODEWRD_IN_q0_0_155;
    rand LDPC_DEC_CODEWRD_IN_q0_0_156_reg_model LDPC_DEC_CODEWRD_IN_q0_0_156;
    rand LDPC_DEC_CODEWRD_IN_q0_0_157_reg_model LDPC_DEC_CODEWRD_IN_q0_0_157;
    rand LDPC_DEC_CODEWRD_IN_q0_0_158_reg_model LDPC_DEC_CODEWRD_IN_q0_0_158;
    rand LDPC_DEC_CODEWRD_IN_q0_0_159_reg_model LDPC_DEC_CODEWRD_IN_q0_0_159;
    rand LDPC_DEC_CODEWRD_IN_q0_0_160_reg_model LDPC_DEC_CODEWRD_IN_q0_0_160;
    rand LDPC_DEC_CODEWRD_IN_q0_0_161_reg_model LDPC_DEC_CODEWRD_IN_q0_0_161;
    rand LDPC_DEC_CODEWRD_IN_q0_0_162_reg_model LDPC_DEC_CODEWRD_IN_q0_0_162;
    rand LDPC_DEC_CODEWRD_IN_q0_0_163_reg_model LDPC_DEC_CODEWRD_IN_q0_0_163;
    rand LDPC_DEC_CODEWRD_IN_q0_0_164_reg_model LDPC_DEC_CODEWRD_IN_q0_0_164;
    rand LDPC_DEC_CODEWRD_IN_q0_0_165_reg_model LDPC_DEC_CODEWRD_IN_q0_0_165;
    rand LDPC_DEC_CODEWRD_IN_q0_0_166_reg_model LDPC_DEC_CODEWRD_IN_q0_0_166;
    rand LDPC_DEC_CODEWRD_IN_q0_0_167_reg_model LDPC_DEC_CODEWRD_IN_q0_0_167;
    rand LDPC_DEC_CODEWRD_IN_q0_0_168_reg_model LDPC_DEC_CODEWRD_IN_q0_0_168;
    rand LDPC_DEC_CODEWRD_IN_q0_0_169_reg_model LDPC_DEC_CODEWRD_IN_q0_0_169;
    rand LDPC_DEC_CODEWRD_IN_q0_0_170_reg_model LDPC_DEC_CODEWRD_IN_q0_0_170;
    rand LDPC_DEC_CODEWRD_IN_q0_0_171_reg_model LDPC_DEC_CODEWRD_IN_q0_0_171;
    rand LDPC_DEC_CODEWRD_IN_q0_0_172_reg_model LDPC_DEC_CODEWRD_IN_q0_0_172;
    rand LDPC_DEC_CODEWRD_IN_q0_0_173_reg_model LDPC_DEC_CODEWRD_IN_q0_0_173;
    rand LDPC_DEC_CODEWRD_IN_q0_0_174_reg_model LDPC_DEC_CODEWRD_IN_q0_0_174;
    rand LDPC_DEC_CODEWRD_IN_q0_0_175_reg_model LDPC_DEC_CODEWRD_IN_q0_0_175;
    rand LDPC_DEC_CODEWRD_IN_q0_0_176_reg_model LDPC_DEC_CODEWRD_IN_q0_0_176;
    rand LDPC_DEC_CODEWRD_IN_q0_0_177_reg_model LDPC_DEC_CODEWRD_IN_q0_0_177;
    rand LDPC_DEC_CODEWRD_IN_q0_0_178_reg_model LDPC_DEC_CODEWRD_IN_q0_0_178;
    rand LDPC_DEC_CODEWRD_IN_q0_0_179_reg_model LDPC_DEC_CODEWRD_IN_q0_0_179;
    rand LDPC_DEC_CODEWRD_IN_q0_0_180_reg_model LDPC_DEC_CODEWRD_IN_q0_0_180;
    rand LDPC_DEC_CODEWRD_IN_q0_0_181_reg_model LDPC_DEC_CODEWRD_IN_q0_0_181;
    rand LDPC_DEC_CODEWRD_IN_q0_0_182_reg_model LDPC_DEC_CODEWRD_IN_q0_0_182;
    rand LDPC_DEC_CODEWRD_IN_q0_0_183_reg_model LDPC_DEC_CODEWRD_IN_q0_0_183;
    rand LDPC_DEC_CODEWRD_IN_q0_0_184_reg_model LDPC_DEC_CODEWRD_IN_q0_0_184;
    rand LDPC_DEC_CODEWRD_IN_q0_0_185_reg_model LDPC_DEC_CODEWRD_IN_q0_0_185;
    rand LDPC_DEC_CODEWRD_IN_q0_0_186_reg_model LDPC_DEC_CODEWRD_IN_q0_0_186;
    rand LDPC_DEC_CODEWRD_IN_q0_0_187_reg_model LDPC_DEC_CODEWRD_IN_q0_0_187;
    rand LDPC_DEC_CODEWRD_IN_q0_0_188_reg_model LDPC_DEC_CODEWRD_IN_q0_0_188;
    rand LDPC_DEC_CODEWRD_IN_q0_0_189_reg_model LDPC_DEC_CODEWRD_IN_q0_0_189;
    rand LDPC_DEC_CODEWRD_IN_q0_0_190_reg_model LDPC_DEC_CODEWRD_IN_q0_0_190;
    rand LDPC_DEC_CODEWRD_IN_q0_0_191_reg_model LDPC_DEC_CODEWRD_IN_q0_0_191;
    rand LDPC_DEC_CODEWRD_IN_q0_0_192_reg_model LDPC_DEC_CODEWRD_IN_q0_0_192;
    rand LDPC_DEC_CODEWRD_IN_q0_0_193_reg_model LDPC_DEC_CODEWRD_IN_q0_0_193;
    rand LDPC_DEC_CODEWRD_IN_q0_0_194_reg_model LDPC_DEC_CODEWRD_IN_q0_0_194;
    rand LDPC_DEC_CODEWRD_IN_q0_0_195_reg_model LDPC_DEC_CODEWRD_IN_q0_0_195;
    rand LDPC_DEC_CODEWRD_IN_q0_0_196_reg_model LDPC_DEC_CODEWRD_IN_q0_0_196;
    rand LDPC_DEC_CODEWRD_IN_q0_0_197_reg_model LDPC_DEC_CODEWRD_IN_q0_0_197;
    rand LDPC_DEC_CODEWRD_IN_q0_0_198_reg_model LDPC_DEC_CODEWRD_IN_q0_0_198;
    rand LDPC_DEC_CODEWRD_IN_q0_0_199_reg_model LDPC_DEC_CODEWRD_IN_q0_0_199;
    rand LDPC_DEC_CODEWRD_IN_q0_0_200_reg_model LDPC_DEC_CODEWRD_IN_q0_0_200;
    rand LDPC_DEC_CODEWRD_IN_q0_0_201_reg_model LDPC_DEC_CODEWRD_IN_q0_0_201;
    rand LDPC_DEC_CODEWRD_IN_q0_0_202_reg_model LDPC_DEC_CODEWRD_IN_q0_0_202;
    rand LDPC_DEC_CODEWRD_IN_q0_0_203_reg_model LDPC_DEC_CODEWRD_IN_q0_0_203;
    rand LDPC_DEC_CODEWRD_IN_q0_0_204_reg_model LDPC_DEC_CODEWRD_IN_q0_0_204;
    rand LDPC_DEC_CODEWRD_IN_q0_0_205_reg_model LDPC_DEC_CODEWRD_IN_q0_0_205;
    rand LDPC_DEC_CODEWRD_IN_q0_0_206_reg_model LDPC_DEC_CODEWRD_IN_q0_0_206;
    rand LDPC_DEC_CODEWRD_IN_q0_0_207_reg_model LDPC_DEC_CODEWRD_IN_q0_0_207;
    rand LDPC_DEC_CODEWRD_IN_q0_1_0_reg_model LDPC_DEC_CODEWRD_IN_q0_1_0;
    rand LDPC_DEC_CODEWRD_IN_q0_1_1_reg_model LDPC_DEC_CODEWRD_IN_q0_1_1;
    rand LDPC_DEC_CODEWRD_IN_q0_1_2_reg_model LDPC_DEC_CODEWRD_IN_q0_1_2;
    rand LDPC_DEC_CODEWRD_IN_q0_1_3_reg_model LDPC_DEC_CODEWRD_IN_q0_1_3;
    rand LDPC_DEC_CODEWRD_IN_q0_1_4_reg_model LDPC_DEC_CODEWRD_IN_q0_1_4;
    rand LDPC_DEC_CODEWRD_IN_q0_1_5_reg_model LDPC_DEC_CODEWRD_IN_q0_1_5;
    rand LDPC_DEC_CODEWRD_IN_q0_1_6_reg_model LDPC_DEC_CODEWRD_IN_q0_1_6;
    rand LDPC_DEC_CODEWRD_IN_q0_1_7_reg_model LDPC_DEC_CODEWRD_IN_q0_1_7;
    rand LDPC_DEC_CODEWRD_IN_q0_1_8_reg_model LDPC_DEC_CODEWRD_IN_q0_1_8;
    rand LDPC_DEC_CODEWRD_IN_q0_1_9_reg_model LDPC_DEC_CODEWRD_IN_q0_1_9;
    rand LDPC_DEC_CODEWRD_IN_q0_1_10_reg_model LDPC_DEC_CODEWRD_IN_q0_1_10;
    rand LDPC_DEC_CODEWRD_IN_q0_1_11_reg_model LDPC_DEC_CODEWRD_IN_q0_1_11;
    rand LDPC_DEC_CODEWRD_IN_q0_1_12_reg_model LDPC_DEC_CODEWRD_IN_q0_1_12;
    rand LDPC_DEC_CODEWRD_IN_q0_1_13_reg_model LDPC_DEC_CODEWRD_IN_q0_1_13;
    rand LDPC_DEC_CODEWRD_IN_q0_1_14_reg_model LDPC_DEC_CODEWRD_IN_q0_1_14;
    rand LDPC_DEC_CODEWRD_IN_q0_1_15_reg_model LDPC_DEC_CODEWRD_IN_q0_1_15;
    rand LDPC_DEC_CODEWRD_IN_q0_1_16_reg_model LDPC_DEC_CODEWRD_IN_q0_1_16;
    rand LDPC_DEC_CODEWRD_IN_q0_1_17_reg_model LDPC_DEC_CODEWRD_IN_q0_1_17;
    rand LDPC_DEC_CODEWRD_IN_q0_1_18_reg_model LDPC_DEC_CODEWRD_IN_q0_1_18;
    rand LDPC_DEC_CODEWRD_IN_q0_1_19_reg_model LDPC_DEC_CODEWRD_IN_q0_1_19;
    rand LDPC_DEC_CODEWRD_IN_q0_1_20_reg_model LDPC_DEC_CODEWRD_IN_q0_1_20;
    rand LDPC_DEC_CODEWRD_IN_q0_1_21_reg_model LDPC_DEC_CODEWRD_IN_q0_1_21;
    rand LDPC_DEC_CODEWRD_IN_q0_1_22_reg_model LDPC_DEC_CODEWRD_IN_q0_1_22;
    rand LDPC_DEC_CODEWRD_IN_q0_1_23_reg_model LDPC_DEC_CODEWRD_IN_q0_1_23;
    rand LDPC_DEC_CODEWRD_IN_q0_1_24_reg_model LDPC_DEC_CODEWRD_IN_q0_1_24;
    rand LDPC_DEC_CODEWRD_IN_q0_1_25_reg_model LDPC_DEC_CODEWRD_IN_q0_1_25;
    rand LDPC_DEC_CODEWRD_IN_q0_1_26_reg_model LDPC_DEC_CODEWRD_IN_q0_1_26;
    rand LDPC_DEC_CODEWRD_IN_q0_1_27_reg_model LDPC_DEC_CODEWRD_IN_q0_1_27;
    rand LDPC_DEC_CODEWRD_IN_q0_1_28_reg_model LDPC_DEC_CODEWRD_IN_q0_1_28;
    rand LDPC_DEC_CODEWRD_IN_q0_1_29_reg_model LDPC_DEC_CODEWRD_IN_q0_1_29;
    rand LDPC_DEC_CODEWRD_IN_q0_1_30_reg_model LDPC_DEC_CODEWRD_IN_q0_1_30;
    rand LDPC_DEC_CODEWRD_IN_q0_1_31_reg_model LDPC_DEC_CODEWRD_IN_q0_1_31;
    rand LDPC_DEC_CODEWRD_IN_q0_1_32_reg_model LDPC_DEC_CODEWRD_IN_q0_1_32;
    rand LDPC_DEC_CODEWRD_IN_q0_1_33_reg_model LDPC_DEC_CODEWRD_IN_q0_1_33;
    rand LDPC_DEC_CODEWRD_IN_q0_1_34_reg_model LDPC_DEC_CODEWRD_IN_q0_1_34;
    rand LDPC_DEC_CODEWRD_IN_q0_1_35_reg_model LDPC_DEC_CODEWRD_IN_q0_1_35;
    rand LDPC_DEC_CODEWRD_IN_q0_1_36_reg_model LDPC_DEC_CODEWRD_IN_q0_1_36;
    rand LDPC_DEC_CODEWRD_IN_q0_1_37_reg_model LDPC_DEC_CODEWRD_IN_q0_1_37;
    rand LDPC_DEC_CODEWRD_IN_q0_1_38_reg_model LDPC_DEC_CODEWRD_IN_q0_1_38;
    rand LDPC_DEC_CODEWRD_IN_q0_1_39_reg_model LDPC_DEC_CODEWRD_IN_q0_1_39;
    rand LDPC_DEC_CODEWRD_IN_q0_1_40_reg_model LDPC_DEC_CODEWRD_IN_q0_1_40;
    rand LDPC_DEC_CODEWRD_IN_q0_1_41_reg_model LDPC_DEC_CODEWRD_IN_q0_1_41;
    rand LDPC_DEC_CODEWRD_IN_q0_1_42_reg_model LDPC_DEC_CODEWRD_IN_q0_1_42;
    rand LDPC_DEC_CODEWRD_IN_q0_1_43_reg_model LDPC_DEC_CODEWRD_IN_q0_1_43;
    rand LDPC_DEC_CODEWRD_IN_q0_1_44_reg_model LDPC_DEC_CODEWRD_IN_q0_1_44;
    rand LDPC_DEC_CODEWRD_IN_q0_1_45_reg_model LDPC_DEC_CODEWRD_IN_q0_1_45;
    rand LDPC_DEC_CODEWRD_IN_q0_1_46_reg_model LDPC_DEC_CODEWRD_IN_q0_1_46;
    rand LDPC_DEC_CODEWRD_IN_q0_1_47_reg_model LDPC_DEC_CODEWRD_IN_q0_1_47;
    rand LDPC_DEC_CODEWRD_IN_q0_1_48_reg_model LDPC_DEC_CODEWRD_IN_q0_1_48;
    rand LDPC_DEC_CODEWRD_IN_q0_1_49_reg_model LDPC_DEC_CODEWRD_IN_q0_1_49;
    rand LDPC_DEC_CODEWRD_IN_q0_1_50_reg_model LDPC_DEC_CODEWRD_IN_q0_1_50;
    rand LDPC_DEC_CODEWRD_IN_q0_1_51_reg_model LDPC_DEC_CODEWRD_IN_q0_1_51;
    rand LDPC_DEC_CODEWRD_IN_q0_1_52_reg_model LDPC_DEC_CODEWRD_IN_q0_1_52;
    rand LDPC_DEC_CODEWRD_IN_q0_1_53_reg_model LDPC_DEC_CODEWRD_IN_q0_1_53;
    rand LDPC_DEC_CODEWRD_IN_q0_1_54_reg_model LDPC_DEC_CODEWRD_IN_q0_1_54;
    rand LDPC_DEC_CODEWRD_IN_q0_1_55_reg_model LDPC_DEC_CODEWRD_IN_q0_1_55;
    rand LDPC_DEC_CODEWRD_IN_q0_1_56_reg_model LDPC_DEC_CODEWRD_IN_q0_1_56;
    rand LDPC_DEC_CODEWRD_IN_q0_1_57_reg_model LDPC_DEC_CODEWRD_IN_q0_1_57;
    rand LDPC_DEC_CODEWRD_IN_q0_1_58_reg_model LDPC_DEC_CODEWRD_IN_q0_1_58;
    rand LDPC_DEC_CODEWRD_IN_q0_1_59_reg_model LDPC_DEC_CODEWRD_IN_q0_1_59;
    rand LDPC_DEC_CODEWRD_IN_q0_1_60_reg_model LDPC_DEC_CODEWRD_IN_q0_1_60;
    rand LDPC_DEC_CODEWRD_IN_q0_1_61_reg_model LDPC_DEC_CODEWRD_IN_q0_1_61;
    rand LDPC_DEC_CODEWRD_IN_q0_1_62_reg_model LDPC_DEC_CODEWRD_IN_q0_1_62;
    rand LDPC_DEC_CODEWRD_IN_q0_1_63_reg_model LDPC_DEC_CODEWRD_IN_q0_1_63;
    rand LDPC_DEC_CODEWRD_IN_q0_1_64_reg_model LDPC_DEC_CODEWRD_IN_q0_1_64;
    rand LDPC_DEC_CODEWRD_IN_q0_1_65_reg_model LDPC_DEC_CODEWRD_IN_q0_1_65;
    rand LDPC_DEC_CODEWRD_IN_q0_1_66_reg_model LDPC_DEC_CODEWRD_IN_q0_1_66;
    rand LDPC_DEC_CODEWRD_IN_q0_1_67_reg_model LDPC_DEC_CODEWRD_IN_q0_1_67;
    rand LDPC_DEC_CODEWRD_IN_q0_1_68_reg_model LDPC_DEC_CODEWRD_IN_q0_1_68;
    rand LDPC_DEC_CODEWRD_IN_q0_1_69_reg_model LDPC_DEC_CODEWRD_IN_q0_1_69;
    rand LDPC_DEC_CODEWRD_IN_q0_1_70_reg_model LDPC_DEC_CODEWRD_IN_q0_1_70;
    rand LDPC_DEC_CODEWRD_IN_q0_1_71_reg_model LDPC_DEC_CODEWRD_IN_q0_1_71;
    rand LDPC_DEC_CODEWRD_IN_q0_1_72_reg_model LDPC_DEC_CODEWRD_IN_q0_1_72;
    rand LDPC_DEC_CODEWRD_IN_q0_1_73_reg_model LDPC_DEC_CODEWRD_IN_q0_1_73;
    rand LDPC_DEC_CODEWRD_IN_q0_1_74_reg_model LDPC_DEC_CODEWRD_IN_q0_1_74;
    rand LDPC_DEC_CODEWRD_IN_q0_1_75_reg_model LDPC_DEC_CODEWRD_IN_q0_1_75;
    rand LDPC_DEC_CODEWRD_IN_q0_1_76_reg_model LDPC_DEC_CODEWRD_IN_q0_1_76;
    rand LDPC_DEC_CODEWRD_IN_q0_1_77_reg_model LDPC_DEC_CODEWRD_IN_q0_1_77;
    rand LDPC_DEC_CODEWRD_IN_q0_1_78_reg_model LDPC_DEC_CODEWRD_IN_q0_1_78;
    rand LDPC_DEC_CODEWRD_IN_q0_1_79_reg_model LDPC_DEC_CODEWRD_IN_q0_1_79;
    rand LDPC_DEC_CODEWRD_IN_q0_1_80_reg_model LDPC_DEC_CODEWRD_IN_q0_1_80;
    rand LDPC_DEC_CODEWRD_IN_q0_1_81_reg_model LDPC_DEC_CODEWRD_IN_q0_1_81;
    rand LDPC_DEC_CODEWRD_IN_q0_1_82_reg_model LDPC_DEC_CODEWRD_IN_q0_1_82;
    rand LDPC_DEC_CODEWRD_IN_q0_1_83_reg_model LDPC_DEC_CODEWRD_IN_q0_1_83;
    rand LDPC_DEC_CODEWRD_IN_q0_1_84_reg_model LDPC_DEC_CODEWRD_IN_q0_1_84;
    rand LDPC_DEC_CODEWRD_IN_q0_1_85_reg_model LDPC_DEC_CODEWRD_IN_q0_1_85;
    rand LDPC_DEC_CODEWRD_IN_q0_1_86_reg_model LDPC_DEC_CODEWRD_IN_q0_1_86;
    rand LDPC_DEC_CODEWRD_IN_q0_1_87_reg_model LDPC_DEC_CODEWRD_IN_q0_1_87;
    rand LDPC_DEC_CODEWRD_IN_q0_1_88_reg_model LDPC_DEC_CODEWRD_IN_q0_1_88;
    rand LDPC_DEC_CODEWRD_IN_q0_1_89_reg_model LDPC_DEC_CODEWRD_IN_q0_1_89;
    rand LDPC_DEC_CODEWRD_IN_q0_1_90_reg_model LDPC_DEC_CODEWRD_IN_q0_1_90;
    rand LDPC_DEC_CODEWRD_IN_q0_1_91_reg_model LDPC_DEC_CODEWRD_IN_q0_1_91;
    rand LDPC_DEC_CODEWRD_IN_q0_1_92_reg_model LDPC_DEC_CODEWRD_IN_q0_1_92;
    rand LDPC_DEC_CODEWRD_IN_q0_1_93_reg_model LDPC_DEC_CODEWRD_IN_q0_1_93;
    rand LDPC_DEC_CODEWRD_IN_q0_1_94_reg_model LDPC_DEC_CODEWRD_IN_q0_1_94;
    rand LDPC_DEC_CODEWRD_IN_q0_1_95_reg_model LDPC_DEC_CODEWRD_IN_q0_1_95;
    rand LDPC_DEC_CODEWRD_IN_q0_1_96_reg_model LDPC_DEC_CODEWRD_IN_q0_1_96;
    rand LDPC_DEC_CODEWRD_IN_q0_1_97_reg_model LDPC_DEC_CODEWRD_IN_q0_1_97;
    rand LDPC_DEC_CODEWRD_IN_q0_1_98_reg_model LDPC_DEC_CODEWRD_IN_q0_1_98;
    rand LDPC_DEC_CODEWRD_IN_q0_1_99_reg_model LDPC_DEC_CODEWRD_IN_q0_1_99;
    rand LDPC_DEC_CODEWRD_IN_q0_1_100_reg_model LDPC_DEC_CODEWRD_IN_q0_1_100;
    rand LDPC_DEC_CODEWRD_IN_q0_1_101_reg_model LDPC_DEC_CODEWRD_IN_q0_1_101;
    rand LDPC_DEC_CODEWRD_IN_q0_1_102_reg_model LDPC_DEC_CODEWRD_IN_q0_1_102;
    rand LDPC_DEC_CODEWRD_IN_q0_1_103_reg_model LDPC_DEC_CODEWRD_IN_q0_1_103;
    rand LDPC_DEC_CODEWRD_IN_q0_1_104_reg_model LDPC_DEC_CODEWRD_IN_q0_1_104;
    rand LDPC_DEC_CODEWRD_IN_q0_1_105_reg_model LDPC_DEC_CODEWRD_IN_q0_1_105;
    rand LDPC_DEC_CODEWRD_IN_q0_1_106_reg_model LDPC_DEC_CODEWRD_IN_q0_1_106;
    rand LDPC_DEC_CODEWRD_IN_q0_1_107_reg_model LDPC_DEC_CODEWRD_IN_q0_1_107;
    rand LDPC_DEC_CODEWRD_IN_q0_1_108_reg_model LDPC_DEC_CODEWRD_IN_q0_1_108;
    rand LDPC_DEC_CODEWRD_IN_q0_1_109_reg_model LDPC_DEC_CODEWRD_IN_q0_1_109;
    rand LDPC_DEC_CODEWRD_IN_q0_1_110_reg_model LDPC_DEC_CODEWRD_IN_q0_1_110;
    rand LDPC_DEC_CODEWRD_IN_q0_1_111_reg_model LDPC_DEC_CODEWRD_IN_q0_1_111;
    rand LDPC_DEC_CODEWRD_IN_q0_1_112_reg_model LDPC_DEC_CODEWRD_IN_q0_1_112;
    rand LDPC_DEC_CODEWRD_IN_q0_1_113_reg_model LDPC_DEC_CODEWRD_IN_q0_1_113;
    rand LDPC_DEC_CODEWRD_IN_q0_1_114_reg_model LDPC_DEC_CODEWRD_IN_q0_1_114;
    rand LDPC_DEC_CODEWRD_IN_q0_1_115_reg_model LDPC_DEC_CODEWRD_IN_q0_1_115;
    rand LDPC_DEC_CODEWRD_IN_q0_1_116_reg_model LDPC_DEC_CODEWRD_IN_q0_1_116;
    rand LDPC_DEC_CODEWRD_IN_q0_1_117_reg_model LDPC_DEC_CODEWRD_IN_q0_1_117;
    rand LDPC_DEC_CODEWRD_IN_q0_1_118_reg_model LDPC_DEC_CODEWRD_IN_q0_1_118;
    rand LDPC_DEC_CODEWRD_IN_q0_1_119_reg_model LDPC_DEC_CODEWRD_IN_q0_1_119;
    rand LDPC_DEC_CODEWRD_IN_q0_1_120_reg_model LDPC_DEC_CODEWRD_IN_q0_1_120;
    rand LDPC_DEC_CODEWRD_IN_q0_1_121_reg_model LDPC_DEC_CODEWRD_IN_q0_1_121;
    rand LDPC_DEC_CODEWRD_IN_q0_1_122_reg_model LDPC_DEC_CODEWRD_IN_q0_1_122;
    rand LDPC_DEC_CODEWRD_IN_q0_1_123_reg_model LDPC_DEC_CODEWRD_IN_q0_1_123;
    rand LDPC_DEC_CODEWRD_IN_q0_1_124_reg_model LDPC_DEC_CODEWRD_IN_q0_1_124;
    rand LDPC_DEC_CODEWRD_IN_q0_1_125_reg_model LDPC_DEC_CODEWRD_IN_q0_1_125;
    rand LDPC_DEC_CODEWRD_IN_q0_1_126_reg_model LDPC_DEC_CODEWRD_IN_q0_1_126;
    rand LDPC_DEC_CODEWRD_IN_q0_1_127_reg_model LDPC_DEC_CODEWRD_IN_q0_1_127;
    rand LDPC_DEC_CODEWRD_IN_q0_1_128_reg_model LDPC_DEC_CODEWRD_IN_q0_1_128;
    rand LDPC_DEC_CODEWRD_IN_q0_1_129_reg_model LDPC_DEC_CODEWRD_IN_q0_1_129;
    rand LDPC_DEC_CODEWRD_IN_q0_1_130_reg_model LDPC_DEC_CODEWRD_IN_q0_1_130;
    rand LDPC_DEC_CODEWRD_IN_q0_1_131_reg_model LDPC_DEC_CODEWRD_IN_q0_1_131;
    rand LDPC_DEC_CODEWRD_IN_q0_1_132_reg_model LDPC_DEC_CODEWRD_IN_q0_1_132;
    rand LDPC_DEC_CODEWRD_IN_q0_1_133_reg_model LDPC_DEC_CODEWRD_IN_q0_1_133;
    rand LDPC_DEC_CODEWRD_IN_q0_1_134_reg_model LDPC_DEC_CODEWRD_IN_q0_1_134;
    rand LDPC_DEC_CODEWRD_IN_q0_1_135_reg_model LDPC_DEC_CODEWRD_IN_q0_1_135;
    rand LDPC_DEC_CODEWRD_IN_q0_1_136_reg_model LDPC_DEC_CODEWRD_IN_q0_1_136;
    rand LDPC_DEC_CODEWRD_IN_q0_1_137_reg_model LDPC_DEC_CODEWRD_IN_q0_1_137;
    rand LDPC_DEC_CODEWRD_IN_q0_1_138_reg_model LDPC_DEC_CODEWRD_IN_q0_1_138;
    rand LDPC_DEC_CODEWRD_IN_q0_1_139_reg_model LDPC_DEC_CODEWRD_IN_q0_1_139;
    rand LDPC_DEC_CODEWRD_IN_q0_1_140_reg_model LDPC_DEC_CODEWRD_IN_q0_1_140;
    rand LDPC_DEC_CODEWRD_IN_q0_1_141_reg_model LDPC_DEC_CODEWRD_IN_q0_1_141;
    rand LDPC_DEC_CODEWRD_IN_q0_1_142_reg_model LDPC_DEC_CODEWRD_IN_q0_1_142;
    rand LDPC_DEC_CODEWRD_IN_q0_1_143_reg_model LDPC_DEC_CODEWRD_IN_q0_1_143;
    rand LDPC_DEC_CODEWRD_IN_q0_1_144_reg_model LDPC_DEC_CODEWRD_IN_q0_1_144;
    rand LDPC_DEC_CODEWRD_IN_q0_1_145_reg_model LDPC_DEC_CODEWRD_IN_q0_1_145;
    rand LDPC_DEC_CODEWRD_IN_q0_1_146_reg_model LDPC_DEC_CODEWRD_IN_q0_1_146;
    rand LDPC_DEC_CODEWRD_IN_q0_1_147_reg_model LDPC_DEC_CODEWRD_IN_q0_1_147;
    rand LDPC_DEC_CODEWRD_IN_q0_1_148_reg_model LDPC_DEC_CODEWRD_IN_q0_1_148;
    rand LDPC_DEC_CODEWRD_IN_q0_1_149_reg_model LDPC_DEC_CODEWRD_IN_q0_1_149;
    rand LDPC_DEC_CODEWRD_IN_q0_1_150_reg_model LDPC_DEC_CODEWRD_IN_q0_1_150;
    rand LDPC_DEC_CODEWRD_IN_q0_1_151_reg_model LDPC_DEC_CODEWRD_IN_q0_1_151;
    rand LDPC_DEC_CODEWRD_IN_q0_1_152_reg_model LDPC_DEC_CODEWRD_IN_q0_1_152;
    rand LDPC_DEC_CODEWRD_IN_q0_1_153_reg_model LDPC_DEC_CODEWRD_IN_q0_1_153;
    rand LDPC_DEC_CODEWRD_IN_q0_1_154_reg_model LDPC_DEC_CODEWRD_IN_q0_1_154;
    rand LDPC_DEC_CODEWRD_IN_q0_1_155_reg_model LDPC_DEC_CODEWRD_IN_q0_1_155;
    rand LDPC_DEC_CODEWRD_IN_q0_1_156_reg_model LDPC_DEC_CODEWRD_IN_q0_1_156;
    rand LDPC_DEC_CODEWRD_IN_q0_1_157_reg_model LDPC_DEC_CODEWRD_IN_q0_1_157;
    rand LDPC_DEC_CODEWRD_IN_q0_1_158_reg_model LDPC_DEC_CODEWRD_IN_q0_1_158;
    rand LDPC_DEC_CODEWRD_IN_q0_1_159_reg_model LDPC_DEC_CODEWRD_IN_q0_1_159;
    rand LDPC_DEC_CODEWRD_IN_q0_1_160_reg_model LDPC_DEC_CODEWRD_IN_q0_1_160;
    rand LDPC_DEC_CODEWRD_IN_q0_1_161_reg_model LDPC_DEC_CODEWRD_IN_q0_1_161;
    rand LDPC_DEC_CODEWRD_IN_q0_1_162_reg_model LDPC_DEC_CODEWRD_IN_q0_1_162;
    rand LDPC_DEC_CODEWRD_IN_q0_1_163_reg_model LDPC_DEC_CODEWRD_IN_q0_1_163;
    rand LDPC_DEC_CODEWRD_IN_q0_1_164_reg_model LDPC_DEC_CODEWRD_IN_q0_1_164;
    rand LDPC_DEC_CODEWRD_IN_q0_1_165_reg_model LDPC_DEC_CODEWRD_IN_q0_1_165;
    rand LDPC_DEC_CODEWRD_IN_q0_1_166_reg_model LDPC_DEC_CODEWRD_IN_q0_1_166;
    rand LDPC_DEC_CODEWRD_IN_q0_1_167_reg_model LDPC_DEC_CODEWRD_IN_q0_1_167;
    rand LDPC_DEC_CODEWRD_IN_q0_1_168_reg_model LDPC_DEC_CODEWRD_IN_q0_1_168;
    rand LDPC_DEC_CODEWRD_IN_q0_1_169_reg_model LDPC_DEC_CODEWRD_IN_q0_1_169;
    rand LDPC_DEC_CODEWRD_IN_q0_1_170_reg_model LDPC_DEC_CODEWRD_IN_q0_1_170;
    rand LDPC_DEC_CODEWRD_IN_q0_1_171_reg_model LDPC_DEC_CODEWRD_IN_q0_1_171;
    rand LDPC_DEC_CODEWRD_IN_q0_1_172_reg_model LDPC_DEC_CODEWRD_IN_q0_1_172;
    rand LDPC_DEC_CODEWRD_IN_q0_1_173_reg_model LDPC_DEC_CODEWRD_IN_q0_1_173;
    rand LDPC_DEC_CODEWRD_IN_q0_1_174_reg_model LDPC_DEC_CODEWRD_IN_q0_1_174;
    rand LDPC_DEC_CODEWRD_IN_q0_1_175_reg_model LDPC_DEC_CODEWRD_IN_q0_1_175;
    rand LDPC_DEC_CODEWRD_IN_q0_1_176_reg_model LDPC_DEC_CODEWRD_IN_q0_1_176;
    rand LDPC_DEC_CODEWRD_IN_q0_1_177_reg_model LDPC_DEC_CODEWRD_IN_q0_1_177;
    rand LDPC_DEC_CODEWRD_IN_q0_1_178_reg_model LDPC_DEC_CODEWRD_IN_q0_1_178;
    rand LDPC_DEC_CODEWRD_IN_q0_1_179_reg_model LDPC_DEC_CODEWRD_IN_q0_1_179;
    rand LDPC_DEC_CODEWRD_IN_q0_1_180_reg_model LDPC_DEC_CODEWRD_IN_q0_1_180;
    rand LDPC_DEC_CODEWRD_IN_q0_1_181_reg_model LDPC_DEC_CODEWRD_IN_q0_1_181;
    rand LDPC_DEC_CODEWRD_IN_q0_1_182_reg_model LDPC_DEC_CODEWRD_IN_q0_1_182;
    rand LDPC_DEC_CODEWRD_IN_q0_1_183_reg_model LDPC_DEC_CODEWRD_IN_q0_1_183;
    rand LDPC_DEC_CODEWRD_IN_q0_1_184_reg_model LDPC_DEC_CODEWRD_IN_q0_1_184;
    rand LDPC_DEC_CODEWRD_IN_q0_1_185_reg_model LDPC_DEC_CODEWRD_IN_q0_1_185;
    rand LDPC_DEC_CODEWRD_IN_q0_1_186_reg_model LDPC_DEC_CODEWRD_IN_q0_1_186;
    rand LDPC_DEC_CODEWRD_IN_q0_1_187_reg_model LDPC_DEC_CODEWRD_IN_q0_1_187;
    rand LDPC_DEC_CODEWRD_IN_q0_1_188_reg_model LDPC_DEC_CODEWRD_IN_q0_1_188;
    rand LDPC_DEC_CODEWRD_IN_q0_1_189_reg_model LDPC_DEC_CODEWRD_IN_q0_1_189;
    rand LDPC_DEC_CODEWRD_IN_q0_1_190_reg_model LDPC_DEC_CODEWRD_IN_q0_1_190;
    rand LDPC_DEC_CODEWRD_IN_q0_1_191_reg_model LDPC_DEC_CODEWRD_IN_q0_1_191;
    rand LDPC_DEC_CODEWRD_IN_q0_1_192_reg_model LDPC_DEC_CODEWRD_IN_q0_1_192;
    rand LDPC_DEC_CODEWRD_IN_q0_1_193_reg_model LDPC_DEC_CODEWRD_IN_q0_1_193;
    rand LDPC_DEC_CODEWRD_IN_q0_1_194_reg_model LDPC_DEC_CODEWRD_IN_q0_1_194;
    rand LDPC_DEC_CODEWRD_IN_q0_1_195_reg_model LDPC_DEC_CODEWRD_IN_q0_1_195;
    rand LDPC_DEC_CODEWRD_IN_q0_1_196_reg_model LDPC_DEC_CODEWRD_IN_q0_1_196;
    rand LDPC_DEC_CODEWRD_IN_q0_1_197_reg_model LDPC_DEC_CODEWRD_IN_q0_1_197;
    rand LDPC_DEC_CODEWRD_IN_q0_1_198_reg_model LDPC_DEC_CODEWRD_IN_q0_1_198;
    rand LDPC_DEC_CODEWRD_IN_q0_1_199_reg_model LDPC_DEC_CODEWRD_IN_q0_1_199;
    rand LDPC_DEC_CODEWRD_IN_q0_1_200_reg_model LDPC_DEC_CODEWRD_IN_q0_1_200;
    rand LDPC_DEC_CODEWRD_IN_q0_1_201_reg_model LDPC_DEC_CODEWRD_IN_q0_1_201;
    rand LDPC_DEC_CODEWRD_IN_q0_1_202_reg_model LDPC_DEC_CODEWRD_IN_q0_1_202;
    rand LDPC_DEC_CODEWRD_IN_q0_1_203_reg_model LDPC_DEC_CODEWRD_IN_q0_1_203;
    rand LDPC_DEC_CODEWRD_IN_q0_1_204_reg_model LDPC_DEC_CODEWRD_IN_q0_1_204;
    rand LDPC_DEC_CODEWRD_IN_q0_1_205_reg_model LDPC_DEC_CODEWRD_IN_q0_1_205;
    rand LDPC_DEC_CODEWRD_IN_q0_1_206_reg_model LDPC_DEC_CODEWRD_IN_q0_1_206;
    rand LDPC_DEC_CODEWRD_IN_q0_1_207_reg_model LDPC_DEC_CODEWRD_IN_q0_1_207;
    rand LDPC_DEC_err_intro_decoder_reg_model LDPC_DEC_err_intro_decoder;
    rand LDPC_DEC_EXPSYND_0_reg_model LDPC_DEC_EXPSYND_0;
    rand LDPC_DEC_EXPSYND_1_reg_model LDPC_DEC_EXPSYND_1;
    rand LDPC_DEC_EXPSYND_2_reg_model LDPC_DEC_EXPSYND_2;
    rand LDPC_DEC_EXPSYND_3_reg_model LDPC_DEC_EXPSYND_3;
    rand LDPC_DEC_EXPSYND_4_reg_model LDPC_DEC_EXPSYND_4;
    rand LDPC_DEC_EXPSYND_5_reg_model LDPC_DEC_EXPSYND_5;
    rand LDPC_DEC_EXPSYND_6_reg_model LDPC_DEC_EXPSYND_6;
    rand LDPC_DEC_EXPSYND_7_reg_model LDPC_DEC_EXPSYND_7;
    rand LDPC_DEC_EXPSYND_8_reg_model LDPC_DEC_EXPSYND_8;
    rand LDPC_DEC_EXPSYND_9_reg_model LDPC_DEC_EXPSYND_9;
    rand LDPC_DEC_EXPSYND_10_reg_model LDPC_DEC_EXPSYND_10;
    rand LDPC_DEC_EXPSYND_11_reg_model LDPC_DEC_EXPSYND_11;
    rand LDPC_DEC_EXPSYND_12_reg_model LDPC_DEC_EXPSYND_12;
    rand LDPC_DEC_EXPSYND_13_reg_model LDPC_DEC_EXPSYND_13;
    rand LDPC_DEC_EXPSYND_14_reg_model LDPC_DEC_EXPSYND_14;
    rand LDPC_DEC_EXPSYND_15_reg_model LDPC_DEC_EXPSYND_15;
    rand LDPC_DEC_EXPSYND_16_reg_model LDPC_DEC_EXPSYND_16;
    rand LDPC_DEC_EXPSYND_17_reg_model LDPC_DEC_EXPSYND_17;
    rand LDPC_DEC_EXPSYND_18_reg_model LDPC_DEC_EXPSYND_18;
    rand LDPC_DEC_EXPSYND_19_reg_model LDPC_DEC_EXPSYND_19;
    rand LDPC_DEC_EXPSYND_20_reg_model LDPC_DEC_EXPSYND_20;
    rand LDPC_DEC_EXPSYND_21_reg_model LDPC_DEC_EXPSYND_21;
    rand LDPC_DEC_EXPSYND_22_reg_model LDPC_DEC_EXPSYND_22;
    rand LDPC_DEC_EXPSYND_23_reg_model LDPC_DEC_EXPSYND_23;
    rand LDPC_DEC_EXPSYND_24_reg_model LDPC_DEC_EXPSYND_24;
    rand LDPC_DEC_EXPSYND_25_reg_model LDPC_DEC_EXPSYND_25;
    rand LDPC_DEC_EXPSYND_26_reg_model LDPC_DEC_EXPSYND_26;
    rand LDPC_DEC_EXPSYND_27_reg_model LDPC_DEC_EXPSYND_27;
    rand LDPC_DEC_EXPSYND_28_reg_model LDPC_DEC_EXPSYND_28;
    rand LDPC_DEC_EXPSYND_29_reg_model LDPC_DEC_EXPSYND_29;
    rand LDPC_DEC_EXPSYND_30_reg_model LDPC_DEC_EXPSYND_30;
    rand LDPC_DEC_EXPSYND_31_reg_model LDPC_DEC_EXPSYND_31;
    rand LDPC_DEC_EXPSYND_32_reg_model LDPC_DEC_EXPSYND_32;
    rand LDPC_DEC_EXPSYND_33_reg_model LDPC_DEC_EXPSYND_33;
    rand LDPC_DEC_EXPSYND_34_reg_model LDPC_DEC_EXPSYND_34;
    rand LDPC_DEC_EXPSYND_35_reg_model LDPC_DEC_EXPSYND_35;
    rand LDPC_DEC_EXPSYND_36_reg_model LDPC_DEC_EXPSYND_36;
    rand LDPC_DEC_EXPSYND_37_reg_model LDPC_DEC_EXPSYND_37;
    rand LDPC_DEC_EXPSYND_38_reg_model LDPC_DEC_EXPSYND_38;
    rand LDPC_DEC_EXPSYND_39_reg_model LDPC_DEC_EXPSYND_39;
    rand LDPC_DEC_EXPSYND_40_reg_model LDPC_DEC_EXPSYND_40;
    rand LDPC_DEC_EXPSYND_41_reg_model LDPC_DEC_EXPSYND_41;
    rand LDPC_DEC_EXPSYND_42_reg_model LDPC_DEC_EXPSYND_42;
    rand LDPC_DEC_EXPSYND_43_reg_model LDPC_DEC_EXPSYND_43;
    rand LDPC_DEC_EXPSYND_44_reg_model LDPC_DEC_EXPSYND_44;
    rand LDPC_DEC_EXPSYND_45_reg_model LDPC_DEC_EXPSYND_45;
    rand LDPC_DEC_EXPSYND_46_reg_model LDPC_DEC_EXPSYND_46;
    rand LDPC_DEC_EXPSYND_47_reg_model LDPC_DEC_EXPSYND_47;
    rand LDPC_DEC_EXPSYND_48_reg_model LDPC_DEC_EXPSYND_48;
    rand LDPC_DEC_EXPSYND_49_reg_model LDPC_DEC_EXPSYND_49;
    rand LDPC_DEC_EXPSYND_50_reg_model LDPC_DEC_EXPSYND_50;
    rand LDPC_DEC_EXPSYND_51_reg_model LDPC_DEC_EXPSYND_51;
    rand LDPC_DEC_EXPSYND_52_reg_model LDPC_DEC_EXPSYND_52;
    rand LDPC_DEC_EXPSYND_53_reg_model LDPC_DEC_EXPSYND_53;
    rand LDPC_DEC_EXPSYND_54_reg_model LDPC_DEC_EXPSYND_54;
    rand LDPC_DEC_EXPSYND_55_reg_model LDPC_DEC_EXPSYND_55;
    rand LDPC_DEC_EXPSYND_56_reg_model LDPC_DEC_EXPSYND_56;
    rand LDPC_DEC_EXPSYND_57_reg_model LDPC_DEC_EXPSYND_57;
    rand LDPC_DEC_EXPSYND_58_reg_model LDPC_DEC_EXPSYND_58;
    rand LDPC_DEC_EXPSYND_59_reg_model LDPC_DEC_EXPSYND_59;
    rand LDPC_DEC_EXPSYND_60_reg_model LDPC_DEC_EXPSYND_60;
    rand LDPC_DEC_EXPSYND_61_reg_model LDPC_DEC_EXPSYND_61;
    rand LDPC_DEC_EXPSYND_62_reg_model LDPC_DEC_EXPSYND_62;
    rand LDPC_DEC_EXPSYND_63_reg_model LDPC_DEC_EXPSYND_63;
    rand LDPC_DEC_EXPSYND_64_reg_model LDPC_DEC_EXPSYND_64;
    rand LDPC_DEC_EXPSYND_65_reg_model LDPC_DEC_EXPSYND_65;
    rand LDPC_DEC_EXPSYND_66_reg_model LDPC_DEC_EXPSYND_66;
    rand LDPC_DEC_EXPSYND_67_reg_model LDPC_DEC_EXPSYND_67;
    rand LDPC_DEC_EXPSYND_68_reg_model LDPC_DEC_EXPSYND_68;
    rand LDPC_DEC_EXPSYND_69_reg_model LDPC_DEC_EXPSYND_69;
    rand LDPC_DEC_EXPSYND_70_reg_model LDPC_DEC_EXPSYND_70;
    rand LDPC_DEC_EXPSYND_71_reg_model LDPC_DEC_EXPSYND_71;
    rand LDPC_DEC_EXPSYND_72_reg_model LDPC_DEC_EXPSYND_72;
    rand LDPC_DEC_EXPSYND_73_reg_model LDPC_DEC_EXPSYND_73;
    rand LDPC_DEC_EXPSYND_74_reg_model LDPC_DEC_EXPSYND_74;
    rand LDPC_DEC_EXPSYND_75_reg_model LDPC_DEC_EXPSYND_75;
    rand LDPC_DEC_EXPSYND_76_reg_model LDPC_DEC_EXPSYND_76;
    rand LDPC_DEC_EXPSYND_77_reg_model LDPC_DEC_EXPSYND_77;
    rand LDPC_DEC_EXPSYND_78_reg_model LDPC_DEC_EXPSYND_78;
    rand LDPC_DEC_EXPSYND_79_reg_model LDPC_DEC_EXPSYND_79;
    rand LDPC_DEC_EXPSYND_80_reg_model LDPC_DEC_EXPSYND_80;
    rand LDPC_DEC_EXPSYND_81_reg_model LDPC_DEC_EXPSYND_81;
    rand LDPC_DEC_EXPSYND_82_reg_model LDPC_DEC_EXPSYND_82;
    rand LDPC_DEC_EXPSYND_83_reg_model LDPC_DEC_EXPSYND_83;
    rand LDPC_DEC_EXPSYND_84_reg_model LDPC_DEC_EXPSYND_84;
    rand LDPC_DEC_EXPSYND_85_reg_model LDPC_DEC_EXPSYND_85;
    rand LDPC_DEC_EXPSYND_86_reg_model LDPC_DEC_EXPSYND_86;
    rand LDPC_DEC_EXPSYND_87_reg_model LDPC_DEC_EXPSYND_87;
    rand LDPC_DEC_EXPSYND_88_reg_model LDPC_DEC_EXPSYND_88;
    rand LDPC_DEC_EXPSYND_89_reg_model LDPC_DEC_EXPSYND_89;
    rand LDPC_DEC_EXPSYND_90_reg_model LDPC_DEC_EXPSYND_90;
    rand LDPC_DEC_EXPSYND_91_reg_model LDPC_DEC_EXPSYND_91;
    rand LDPC_DEC_EXPSYND_92_reg_model LDPC_DEC_EXPSYND_92;
    rand LDPC_DEC_EXPSYND_93_reg_model LDPC_DEC_EXPSYND_93;
    rand LDPC_DEC_EXPSYND_94_reg_model LDPC_DEC_EXPSYND_94;
    rand LDPC_DEC_EXPSYND_95_reg_model LDPC_DEC_EXPSYND_95;
    rand LDPC_DEC_EXPSYND_96_reg_model LDPC_DEC_EXPSYND_96;
    rand LDPC_DEC_EXPSYND_97_reg_model LDPC_DEC_EXPSYND_97;
    rand LDPC_DEC_EXPSYND_98_reg_model LDPC_DEC_EXPSYND_98;
    rand LDPC_DEC_EXPSYND_99_reg_model LDPC_DEC_EXPSYND_99;
    rand LDPC_DEC_EXPSYND_100_reg_model LDPC_DEC_EXPSYND_100;
    rand LDPC_DEC_EXPSYND_101_reg_model LDPC_DEC_EXPSYND_101;
    rand LDPC_DEC_EXPSYND_102_reg_model LDPC_DEC_EXPSYND_102;
    rand LDPC_DEC_EXPSYND_103_reg_model LDPC_DEC_EXPSYND_103;
    rand LDPC_DEC_EXPSYND_104_reg_model LDPC_DEC_EXPSYND_104;
    rand LDPC_DEC_EXPSYND_105_reg_model LDPC_DEC_EXPSYND_105;
    rand LDPC_DEC_EXPSYND_106_reg_model LDPC_DEC_EXPSYND_106;
    rand LDPC_DEC_EXPSYND_107_reg_model LDPC_DEC_EXPSYND_107;
    rand LDPC_DEC_EXPSYND_108_reg_model LDPC_DEC_EXPSYND_108;
    rand LDPC_DEC_EXPSYND_109_reg_model LDPC_DEC_EXPSYND_109;
    rand LDPC_DEC_EXPSYND_110_reg_model LDPC_DEC_EXPSYND_110;
    rand LDPC_DEC_EXPSYND_111_reg_model LDPC_DEC_EXPSYND_111;
    rand LDPC_DEC_EXPSYND_112_reg_model LDPC_DEC_EXPSYND_112;
    rand LDPC_DEC_EXPSYND_113_reg_model LDPC_DEC_EXPSYND_113;
    rand LDPC_DEC_EXPSYND_114_reg_model LDPC_DEC_EXPSYND_114;
    rand LDPC_DEC_EXPSYND_115_reg_model LDPC_DEC_EXPSYND_115;
    rand LDPC_DEC_EXPSYND_116_reg_model LDPC_DEC_EXPSYND_116;
    rand LDPC_DEC_EXPSYND_117_reg_model LDPC_DEC_EXPSYND_117;
    rand LDPC_DEC_EXPSYND_118_reg_model LDPC_DEC_EXPSYND_118;
    rand LDPC_DEC_EXPSYND_119_reg_model LDPC_DEC_EXPSYND_119;
    rand LDPC_DEC_EXPSYND_120_reg_model LDPC_DEC_EXPSYND_120;
    rand LDPC_DEC_EXPSYND_121_reg_model LDPC_DEC_EXPSYND_121;
    rand LDPC_DEC_EXPSYND_122_reg_model LDPC_DEC_EXPSYND_122;
    rand LDPC_DEC_EXPSYND_123_reg_model LDPC_DEC_EXPSYND_123;
    rand LDPC_DEC_EXPSYND_124_reg_model LDPC_DEC_EXPSYND_124;
    rand LDPC_DEC_EXPSYND_125_reg_model LDPC_DEC_EXPSYND_125;
    rand LDPC_DEC_EXPSYND_126_reg_model LDPC_DEC_EXPSYND_126;
    rand LDPC_DEC_EXPSYND_127_reg_model LDPC_DEC_EXPSYND_127;
    rand LDPC_DEC_EXPSYND_128_reg_model LDPC_DEC_EXPSYND_128;
    rand LDPC_DEC_EXPSYND_129_reg_model LDPC_DEC_EXPSYND_129;
    rand LDPC_DEC_EXPSYND_130_reg_model LDPC_DEC_EXPSYND_130;
    rand LDPC_DEC_EXPSYND_131_reg_model LDPC_DEC_EXPSYND_131;
    rand LDPC_DEC_EXPSYND_132_reg_model LDPC_DEC_EXPSYND_132;
    rand LDPC_DEC_EXPSYND_133_reg_model LDPC_DEC_EXPSYND_133;
    rand LDPC_DEC_EXPSYND_134_reg_model LDPC_DEC_EXPSYND_134;
    rand LDPC_DEC_EXPSYND_135_reg_model LDPC_DEC_EXPSYND_135;
    rand LDPC_DEC_EXPSYND_136_reg_model LDPC_DEC_EXPSYND_136;
    rand LDPC_DEC_EXPSYND_137_reg_model LDPC_DEC_EXPSYND_137;
    rand LDPC_DEC_EXPSYND_138_reg_model LDPC_DEC_EXPSYND_138;
    rand LDPC_DEC_EXPSYND_139_reg_model LDPC_DEC_EXPSYND_139;
    rand LDPC_DEC_EXPSYND_140_reg_model LDPC_DEC_EXPSYND_140;
    rand LDPC_DEC_EXPSYND_141_reg_model LDPC_DEC_EXPSYND_141;
    rand LDPC_DEC_EXPSYND_142_reg_model LDPC_DEC_EXPSYND_142;
    rand LDPC_DEC_EXPSYND_143_reg_model LDPC_DEC_EXPSYND_143;
    rand LDPC_DEC_EXPSYND_144_reg_model LDPC_DEC_EXPSYND_144;
    rand LDPC_DEC_EXPSYND_145_reg_model LDPC_DEC_EXPSYND_145;
    rand LDPC_DEC_EXPSYND_146_reg_model LDPC_DEC_EXPSYND_146;
    rand LDPC_DEC_EXPSYND_147_reg_model LDPC_DEC_EXPSYND_147;
    rand LDPC_DEC_EXPSYND_148_reg_model LDPC_DEC_EXPSYND_148;
    rand LDPC_DEC_EXPSYND_149_reg_model LDPC_DEC_EXPSYND_149;
    rand LDPC_DEC_EXPSYND_150_reg_model LDPC_DEC_EXPSYND_150;
    rand LDPC_DEC_EXPSYND_151_reg_model LDPC_DEC_EXPSYND_151;
    rand LDPC_DEC_EXPSYND_152_reg_model LDPC_DEC_EXPSYND_152;
    rand LDPC_DEC_EXPSYND_153_reg_model LDPC_DEC_EXPSYND_153;
    rand LDPC_DEC_EXPSYND_154_reg_model LDPC_DEC_EXPSYND_154;
    rand LDPC_DEC_EXPSYND_155_reg_model LDPC_DEC_EXPSYND_155;
    rand LDPC_DEC_EXPSYND_156_reg_model LDPC_DEC_EXPSYND_156;
    rand LDPC_DEC_EXPSYND_157_reg_model LDPC_DEC_EXPSYND_157;
    rand LDPC_DEC_EXPSYND_158_reg_model LDPC_DEC_EXPSYND_158;
    rand LDPC_DEC_EXPSYND_159_reg_model LDPC_DEC_EXPSYND_159;
    rand LDPC_DEC_EXPSYND_160_reg_model LDPC_DEC_EXPSYND_160;
    rand LDPC_DEC_EXPSYND_161_reg_model LDPC_DEC_EXPSYND_161;
    rand LDPC_DEC_EXPSYND_162_reg_model LDPC_DEC_EXPSYND_162;
    rand LDPC_DEC_EXPSYND_163_reg_model LDPC_DEC_EXPSYND_163;
    rand LDPC_DEC_EXPSYND_164_reg_model LDPC_DEC_EXPSYND_164;
    rand LDPC_DEC_EXPSYND_165_reg_model LDPC_DEC_EXPSYND_165;
    rand LDPC_DEC_EXPSYND_166_reg_model LDPC_DEC_EXPSYND_166;
    rand LDPC_DEC_EXPSYND_167_reg_model LDPC_DEC_EXPSYND_167;
    rand LDPC_DEC_PROBABILITY_reg_model LDPC_DEC_PROBABILITY;
    rand LDPC_DEC_HAMDIST_LOOP_MAX_reg_model LDPC_DEC_HAMDIST_LOOP_MAX;
    rand LDPC_DEC_HAMDIST_LOOP_PERCENTAGE_reg_model LDPC_DEC_HAMDIST_LOOP_PERCENTAGE;
    rand LDPC_DEC_HAMDIST_IIR1_reg_model LDPC_DEC_HAMDIST_IIR1;
    rand LDPC_DEC_HAMDIST_IIR2_NOT_USED_reg_model LDPC_DEC_HAMDIST_IIR2_NOT_USED;
    rand LDPC_DEC_HAMDIST_IIR3_NOT_USED_reg_model LDPC_DEC_HAMDIST_IIR3_NOT_USED;
    rand LDPC_DEC_SYN_VALID_CWORD_DEC_final_reg_model LDPC_DEC_SYN_VALID_CWORD_DEC_final;
    rand LDPC_DEC_START_DEC_reg_model LDPC_DEC_START_DEC;
    rand LDPC_DEC_CONVERGED_LOOPS_ENDED_reg_model LDPC_DEC_CONVERGED_LOOPS_ENDED;
    rand LDPC_DEC_CONVERGED_PASS_FAIL_reg_model LDPC_DEC_CONVERGED_PASS_FAIL;
    rand LDPC_DEC_CODEWRD_OUT_BIT_0_reg_model LDPC_DEC_CODEWRD_OUT_BIT_0;
    rand LDPC_DEC_CODEWRD_OUT_BIT_1_reg_model LDPC_DEC_CODEWRD_OUT_BIT_1;
    rand LDPC_DEC_CODEWRD_OUT_BIT_2_reg_model LDPC_DEC_CODEWRD_OUT_BIT_2;
    rand LDPC_DEC_CODEWRD_OUT_BIT_3_reg_model LDPC_DEC_CODEWRD_OUT_BIT_3;
    rand LDPC_DEC_CODEWRD_OUT_BIT_4_reg_model LDPC_DEC_CODEWRD_OUT_BIT_4;
    rand LDPC_DEC_CODEWRD_OUT_BIT_5_reg_model LDPC_DEC_CODEWRD_OUT_BIT_5;
    rand LDPC_DEC_CODEWRD_OUT_BIT_6_reg_model LDPC_DEC_CODEWRD_OUT_BIT_6;
    rand LDPC_DEC_CODEWRD_OUT_BIT_7_reg_model LDPC_DEC_CODEWRD_OUT_BIT_7;
    rand LDPC_DEC_CODEWRD_OUT_BIT_8_reg_model LDPC_DEC_CODEWRD_OUT_BIT_8;
    rand LDPC_DEC_CODEWRD_OUT_BIT_9_reg_model LDPC_DEC_CODEWRD_OUT_BIT_9;
    rand LDPC_DEC_CODEWRD_OUT_BIT_10_reg_model LDPC_DEC_CODEWRD_OUT_BIT_10;
    rand LDPC_DEC_CODEWRD_OUT_BIT_11_reg_model LDPC_DEC_CODEWRD_OUT_BIT_11;
    rand LDPC_DEC_CODEWRD_OUT_BIT_12_reg_model LDPC_DEC_CODEWRD_OUT_BIT_12;
    rand LDPC_DEC_CODEWRD_OUT_BIT_13_reg_model LDPC_DEC_CODEWRD_OUT_BIT_13;
    rand LDPC_DEC_CODEWRD_OUT_BIT_14_reg_model LDPC_DEC_CODEWRD_OUT_BIT_14;
    rand LDPC_DEC_CODEWRD_OUT_BIT_15_reg_model LDPC_DEC_CODEWRD_OUT_BIT_15;
    rand LDPC_DEC_CODEWRD_OUT_BIT_16_reg_model LDPC_DEC_CODEWRD_OUT_BIT_16;
    rand LDPC_DEC_CODEWRD_OUT_BIT_17_reg_model LDPC_DEC_CODEWRD_OUT_BIT_17;
    rand LDPC_DEC_CODEWRD_OUT_BIT_18_reg_model LDPC_DEC_CODEWRD_OUT_BIT_18;
    rand LDPC_DEC_CODEWRD_OUT_BIT_19_reg_model LDPC_DEC_CODEWRD_OUT_BIT_19;
    rand LDPC_DEC_CODEWRD_OUT_BIT_20_reg_model LDPC_DEC_CODEWRD_OUT_BIT_20;
    rand LDPC_DEC_CODEWRD_OUT_BIT_21_reg_model LDPC_DEC_CODEWRD_OUT_BIT_21;
    rand LDPC_DEC_CODEWRD_OUT_BIT_22_reg_model LDPC_DEC_CODEWRD_OUT_BIT_22;
    rand LDPC_DEC_CODEWRD_OUT_BIT_23_reg_model LDPC_DEC_CODEWRD_OUT_BIT_23;
    rand LDPC_DEC_CODEWRD_OUT_BIT_24_reg_model LDPC_DEC_CODEWRD_OUT_BIT_24;
    rand LDPC_DEC_CODEWRD_OUT_BIT_25_reg_model LDPC_DEC_CODEWRD_OUT_BIT_25;
    rand LDPC_DEC_CODEWRD_OUT_BIT_26_reg_model LDPC_DEC_CODEWRD_OUT_BIT_26;
    rand LDPC_DEC_CODEWRD_OUT_BIT_27_reg_model LDPC_DEC_CODEWRD_OUT_BIT_27;
    rand LDPC_DEC_CODEWRD_OUT_BIT_28_reg_model LDPC_DEC_CODEWRD_OUT_BIT_28;
    rand LDPC_DEC_CODEWRD_OUT_BIT_29_reg_model LDPC_DEC_CODEWRD_OUT_BIT_29;
    rand LDPC_DEC_CODEWRD_OUT_BIT_30_reg_model LDPC_DEC_CODEWRD_OUT_BIT_30;
    rand LDPC_DEC_CODEWRD_OUT_BIT_31_reg_model LDPC_DEC_CODEWRD_OUT_BIT_31;
    rand LDPC_DEC_CODEWRD_OUT_BIT_32_reg_model LDPC_DEC_CODEWRD_OUT_BIT_32;
    rand LDPC_DEC_CODEWRD_OUT_BIT_33_reg_model LDPC_DEC_CODEWRD_OUT_BIT_33;
    rand LDPC_DEC_CODEWRD_OUT_BIT_34_reg_model LDPC_DEC_CODEWRD_OUT_BIT_34;
    rand LDPC_DEC_CODEWRD_OUT_BIT_35_reg_model LDPC_DEC_CODEWRD_OUT_BIT_35;
    rand LDPC_DEC_CODEWRD_OUT_BIT_36_reg_model LDPC_DEC_CODEWRD_OUT_BIT_36;
    rand LDPC_DEC_CODEWRD_OUT_BIT_37_reg_model LDPC_DEC_CODEWRD_OUT_BIT_37;
    rand LDPC_DEC_CODEWRD_OUT_BIT_38_reg_model LDPC_DEC_CODEWRD_OUT_BIT_38;
    rand LDPC_DEC_CODEWRD_OUT_BIT_39_reg_model LDPC_DEC_CODEWRD_OUT_BIT_39;
    rand LDPC_DEC_CODEWRD_OUT_BIT_40_reg_model LDPC_DEC_CODEWRD_OUT_BIT_40;
    rand LDPC_DEC_CODEWRD_OUT_BIT_41_reg_model LDPC_DEC_CODEWRD_OUT_BIT_41;
    rand LDPC_DEC_CODEWRD_OUT_BIT_42_reg_model LDPC_DEC_CODEWRD_OUT_BIT_42;
    rand LDPC_DEC_CODEWRD_OUT_BIT_43_reg_model LDPC_DEC_CODEWRD_OUT_BIT_43;
    rand LDPC_DEC_CODEWRD_OUT_BIT_44_reg_model LDPC_DEC_CODEWRD_OUT_BIT_44;
    rand LDPC_DEC_CODEWRD_OUT_BIT_45_reg_model LDPC_DEC_CODEWRD_OUT_BIT_45;
    rand LDPC_DEC_CODEWRD_OUT_BIT_46_reg_model LDPC_DEC_CODEWRD_OUT_BIT_46;
    rand LDPC_DEC_CODEWRD_OUT_BIT_47_reg_model LDPC_DEC_CODEWRD_OUT_BIT_47;
    rand LDPC_DEC_CODEWRD_OUT_BIT_48_reg_model LDPC_DEC_CODEWRD_OUT_BIT_48;
    rand LDPC_DEC_CODEWRD_OUT_BIT_49_reg_model LDPC_DEC_CODEWRD_OUT_BIT_49;
    rand LDPC_DEC_CODEWRD_OUT_BIT_50_reg_model LDPC_DEC_CODEWRD_OUT_BIT_50;
    rand LDPC_DEC_CODEWRD_OUT_BIT_51_reg_model LDPC_DEC_CODEWRD_OUT_BIT_51;
    rand LDPC_DEC_CODEWRD_OUT_BIT_52_reg_model LDPC_DEC_CODEWRD_OUT_BIT_52;
    rand LDPC_DEC_CODEWRD_OUT_BIT_53_reg_model LDPC_DEC_CODEWRD_OUT_BIT_53;
    rand LDPC_DEC_CODEWRD_OUT_BIT_54_reg_model LDPC_DEC_CODEWRD_OUT_BIT_54;
    rand LDPC_DEC_CODEWRD_OUT_BIT_55_reg_model LDPC_DEC_CODEWRD_OUT_BIT_55;
    rand LDPC_DEC_CODEWRD_OUT_BIT_56_reg_model LDPC_DEC_CODEWRD_OUT_BIT_56;
    rand LDPC_DEC_CODEWRD_OUT_BIT_57_reg_model LDPC_DEC_CODEWRD_OUT_BIT_57;
    rand LDPC_DEC_CODEWRD_OUT_BIT_58_reg_model LDPC_DEC_CODEWRD_OUT_BIT_58;
    rand LDPC_DEC_CODEWRD_OUT_BIT_59_reg_model LDPC_DEC_CODEWRD_OUT_BIT_59;
    rand LDPC_DEC_CODEWRD_OUT_BIT_60_reg_model LDPC_DEC_CODEWRD_OUT_BIT_60;
    rand LDPC_DEC_CODEWRD_OUT_BIT_61_reg_model LDPC_DEC_CODEWRD_OUT_BIT_61;
    rand LDPC_DEC_CODEWRD_OUT_BIT_62_reg_model LDPC_DEC_CODEWRD_OUT_BIT_62;
    rand LDPC_DEC_CODEWRD_OUT_BIT_63_reg_model LDPC_DEC_CODEWRD_OUT_BIT_63;
    rand LDPC_DEC_CODEWRD_OUT_BIT_64_reg_model LDPC_DEC_CODEWRD_OUT_BIT_64;
    rand LDPC_DEC_CODEWRD_OUT_BIT_65_reg_model LDPC_DEC_CODEWRD_OUT_BIT_65;
    rand LDPC_DEC_CODEWRD_OUT_BIT_66_reg_model LDPC_DEC_CODEWRD_OUT_BIT_66;
    rand LDPC_DEC_CODEWRD_OUT_BIT_67_reg_model LDPC_DEC_CODEWRD_OUT_BIT_67;
    rand LDPC_DEC_CODEWRD_OUT_BIT_68_reg_model LDPC_DEC_CODEWRD_OUT_BIT_68;
    rand LDPC_DEC_CODEWRD_OUT_BIT_69_reg_model LDPC_DEC_CODEWRD_OUT_BIT_69;
    rand LDPC_DEC_CODEWRD_OUT_BIT_70_reg_model LDPC_DEC_CODEWRD_OUT_BIT_70;
    rand LDPC_DEC_CODEWRD_OUT_BIT_71_reg_model LDPC_DEC_CODEWRD_OUT_BIT_71;
    rand LDPC_DEC_CODEWRD_OUT_BIT_72_reg_model LDPC_DEC_CODEWRD_OUT_BIT_72;
    rand LDPC_DEC_CODEWRD_OUT_BIT_73_reg_model LDPC_DEC_CODEWRD_OUT_BIT_73;
    rand LDPC_DEC_CODEWRD_OUT_BIT_74_reg_model LDPC_DEC_CODEWRD_OUT_BIT_74;
    rand LDPC_DEC_CODEWRD_OUT_BIT_75_reg_model LDPC_DEC_CODEWRD_OUT_BIT_75;
    rand LDPC_DEC_CODEWRD_OUT_BIT_76_reg_model LDPC_DEC_CODEWRD_OUT_BIT_76;
    rand LDPC_DEC_CODEWRD_OUT_BIT_77_reg_model LDPC_DEC_CODEWRD_OUT_BIT_77;
    rand LDPC_DEC_CODEWRD_OUT_BIT_78_reg_model LDPC_DEC_CODEWRD_OUT_BIT_78;
    rand LDPC_DEC_CODEWRD_OUT_BIT_79_reg_model LDPC_DEC_CODEWRD_OUT_BIT_79;
    rand LDPC_DEC_CODEWRD_OUT_BIT_80_reg_model LDPC_DEC_CODEWRD_OUT_BIT_80;
    rand LDPC_DEC_CODEWRD_OUT_BIT_81_reg_model LDPC_DEC_CODEWRD_OUT_BIT_81;
    rand LDPC_DEC_CODEWRD_OUT_BIT_82_reg_model LDPC_DEC_CODEWRD_OUT_BIT_82;
    rand LDPC_DEC_CODEWRD_OUT_BIT_83_reg_model LDPC_DEC_CODEWRD_OUT_BIT_83;
    rand LDPC_DEC_CODEWRD_OUT_BIT_84_reg_model LDPC_DEC_CODEWRD_OUT_BIT_84;
    rand LDPC_DEC_CODEWRD_OUT_BIT_85_reg_model LDPC_DEC_CODEWRD_OUT_BIT_85;
    rand LDPC_DEC_CODEWRD_OUT_BIT_86_reg_model LDPC_DEC_CODEWRD_OUT_BIT_86;
    rand LDPC_DEC_CODEWRD_OUT_BIT_87_reg_model LDPC_DEC_CODEWRD_OUT_BIT_87;
    rand LDPC_DEC_CODEWRD_OUT_BIT_88_reg_model LDPC_DEC_CODEWRD_OUT_BIT_88;
    rand LDPC_DEC_CODEWRD_OUT_BIT_89_reg_model LDPC_DEC_CODEWRD_OUT_BIT_89;
    rand LDPC_DEC_CODEWRD_OUT_BIT_90_reg_model LDPC_DEC_CODEWRD_OUT_BIT_90;
    rand LDPC_DEC_CODEWRD_OUT_BIT_91_reg_model LDPC_DEC_CODEWRD_OUT_BIT_91;
    rand LDPC_DEC_CODEWRD_OUT_BIT_92_reg_model LDPC_DEC_CODEWRD_OUT_BIT_92;
    rand LDPC_DEC_CODEWRD_OUT_BIT_93_reg_model LDPC_DEC_CODEWRD_OUT_BIT_93;
    rand LDPC_DEC_CODEWRD_OUT_BIT_94_reg_model LDPC_DEC_CODEWRD_OUT_BIT_94;
    rand LDPC_DEC_CODEWRD_OUT_BIT_95_reg_model LDPC_DEC_CODEWRD_OUT_BIT_95;
    rand LDPC_DEC_CODEWRD_OUT_BIT_96_reg_model LDPC_DEC_CODEWRD_OUT_BIT_96;
    rand LDPC_DEC_CODEWRD_OUT_BIT_97_reg_model LDPC_DEC_CODEWRD_OUT_BIT_97;
    rand LDPC_DEC_CODEWRD_OUT_BIT_98_reg_model LDPC_DEC_CODEWRD_OUT_BIT_98;
    rand LDPC_DEC_CODEWRD_OUT_BIT_99_reg_model LDPC_DEC_CODEWRD_OUT_BIT_99;
    rand LDPC_DEC_CODEWRD_OUT_BIT_100_reg_model LDPC_DEC_CODEWRD_OUT_BIT_100;
    rand LDPC_DEC_CODEWRD_OUT_BIT_101_reg_model LDPC_DEC_CODEWRD_OUT_BIT_101;
    rand LDPC_DEC_CODEWRD_OUT_BIT_102_reg_model LDPC_DEC_CODEWRD_OUT_BIT_102;
    rand LDPC_DEC_CODEWRD_OUT_BIT_103_reg_model LDPC_DEC_CODEWRD_OUT_BIT_103;
    rand LDPC_DEC_CODEWRD_OUT_BIT_104_reg_model LDPC_DEC_CODEWRD_OUT_BIT_104;
    rand LDPC_DEC_CODEWRD_OUT_BIT_105_reg_model LDPC_DEC_CODEWRD_OUT_BIT_105;
    rand LDPC_DEC_CODEWRD_OUT_BIT_106_reg_model LDPC_DEC_CODEWRD_OUT_BIT_106;
    rand LDPC_DEC_CODEWRD_OUT_BIT_107_reg_model LDPC_DEC_CODEWRD_OUT_BIT_107;
    rand LDPC_DEC_CODEWRD_OUT_BIT_108_reg_model LDPC_DEC_CODEWRD_OUT_BIT_108;
    rand LDPC_DEC_CODEWRD_OUT_BIT_109_reg_model LDPC_DEC_CODEWRD_OUT_BIT_109;
    rand LDPC_DEC_CODEWRD_OUT_BIT_110_reg_model LDPC_DEC_CODEWRD_OUT_BIT_110;
    rand LDPC_DEC_CODEWRD_OUT_BIT_111_reg_model LDPC_DEC_CODEWRD_OUT_BIT_111;
    rand LDPC_DEC_CODEWRD_OUT_BIT_112_reg_model LDPC_DEC_CODEWRD_OUT_BIT_112;
    rand LDPC_DEC_CODEWRD_OUT_BIT_113_reg_model LDPC_DEC_CODEWRD_OUT_BIT_113;
    rand LDPC_DEC_CODEWRD_OUT_BIT_114_reg_model LDPC_DEC_CODEWRD_OUT_BIT_114;
    rand LDPC_DEC_CODEWRD_OUT_BIT_115_reg_model LDPC_DEC_CODEWRD_OUT_BIT_115;
    rand LDPC_DEC_CODEWRD_OUT_BIT_116_reg_model LDPC_DEC_CODEWRD_OUT_BIT_116;
    rand LDPC_DEC_CODEWRD_OUT_BIT_117_reg_model LDPC_DEC_CODEWRD_OUT_BIT_117;
    rand LDPC_DEC_CODEWRD_OUT_BIT_118_reg_model LDPC_DEC_CODEWRD_OUT_BIT_118;
    rand LDPC_DEC_CODEWRD_OUT_BIT_119_reg_model LDPC_DEC_CODEWRD_OUT_BIT_119;
    rand LDPC_DEC_CODEWRD_OUT_BIT_120_reg_model LDPC_DEC_CODEWRD_OUT_BIT_120;
    rand LDPC_DEC_CODEWRD_OUT_BIT_121_reg_model LDPC_DEC_CODEWRD_OUT_BIT_121;
    rand LDPC_DEC_CODEWRD_OUT_BIT_122_reg_model LDPC_DEC_CODEWRD_OUT_BIT_122;
    rand LDPC_DEC_CODEWRD_OUT_BIT_123_reg_model LDPC_DEC_CODEWRD_OUT_BIT_123;
    rand LDPC_DEC_CODEWRD_OUT_BIT_124_reg_model LDPC_DEC_CODEWRD_OUT_BIT_124;
    rand LDPC_DEC_CODEWRD_OUT_BIT_125_reg_model LDPC_DEC_CODEWRD_OUT_BIT_125;
    rand LDPC_DEC_CODEWRD_OUT_BIT_126_reg_model LDPC_DEC_CODEWRD_OUT_BIT_126;
    rand LDPC_DEC_CODEWRD_OUT_BIT_127_reg_model LDPC_DEC_CODEWRD_OUT_BIT_127;
    rand LDPC_DEC_CODEWRD_OUT_BIT_128_reg_model LDPC_DEC_CODEWRD_OUT_BIT_128;
    rand LDPC_DEC_CODEWRD_OUT_BIT_129_reg_model LDPC_DEC_CODEWRD_OUT_BIT_129;
    rand LDPC_DEC_CODEWRD_OUT_BIT_130_reg_model LDPC_DEC_CODEWRD_OUT_BIT_130;
    rand LDPC_DEC_CODEWRD_OUT_BIT_131_reg_model LDPC_DEC_CODEWRD_OUT_BIT_131;
    rand LDPC_DEC_CODEWRD_OUT_BIT_132_reg_model LDPC_DEC_CODEWRD_OUT_BIT_132;
    rand LDPC_DEC_CODEWRD_OUT_BIT_133_reg_model LDPC_DEC_CODEWRD_OUT_BIT_133;
    rand LDPC_DEC_CODEWRD_OUT_BIT_134_reg_model LDPC_DEC_CODEWRD_OUT_BIT_134;
    rand LDPC_DEC_CODEWRD_OUT_BIT_135_reg_model LDPC_DEC_CODEWRD_OUT_BIT_135;
    rand LDPC_DEC_CODEWRD_OUT_BIT_136_reg_model LDPC_DEC_CODEWRD_OUT_BIT_136;
    rand LDPC_DEC_CODEWRD_OUT_BIT_137_reg_model LDPC_DEC_CODEWRD_OUT_BIT_137;
    rand LDPC_DEC_CODEWRD_OUT_BIT_138_reg_model LDPC_DEC_CODEWRD_OUT_BIT_138;
    rand LDPC_DEC_CODEWRD_OUT_BIT_139_reg_model LDPC_DEC_CODEWRD_OUT_BIT_139;
    rand LDPC_DEC_CODEWRD_OUT_BIT_140_reg_model LDPC_DEC_CODEWRD_OUT_BIT_140;
    rand LDPC_DEC_CODEWRD_OUT_BIT_141_reg_model LDPC_DEC_CODEWRD_OUT_BIT_141;
    rand LDPC_DEC_CODEWRD_OUT_BIT_142_reg_model LDPC_DEC_CODEWRD_OUT_BIT_142;
    rand LDPC_DEC_CODEWRD_OUT_BIT_143_reg_model LDPC_DEC_CODEWRD_OUT_BIT_143;
    rand LDPC_DEC_CODEWRD_OUT_BIT_144_reg_model LDPC_DEC_CODEWRD_OUT_BIT_144;
    rand LDPC_DEC_CODEWRD_OUT_BIT_145_reg_model LDPC_DEC_CODEWRD_OUT_BIT_145;
    rand LDPC_DEC_CODEWRD_OUT_BIT_146_reg_model LDPC_DEC_CODEWRD_OUT_BIT_146;
    rand LDPC_DEC_CODEWRD_OUT_BIT_147_reg_model LDPC_DEC_CODEWRD_OUT_BIT_147;
    rand LDPC_DEC_CODEWRD_OUT_BIT_148_reg_model LDPC_DEC_CODEWRD_OUT_BIT_148;
    rand LDPC_DEC_CODEWRD_OUT_BIT_149_reg_model LDPC_DEC_CODEWRD_OUT_BIT_149;
    rand LDPC_DEC_CODEWRD_OUT_BIT_150_reg_model LDPC_DEC_CODEWRD_OUT_BIT_150;
    rand LDPC_DEC_CODEWRD_OUT_BIT_151_reg_model LDPC_DEC_CODEWRD_OUT_BIT_151;
    rand LDPC_DEC_CODEWRD_OUT_BIT_152_reg_model LDPC_DEC_CODEWRD_OUT_BIT_152;
    rand LDPC_DEC_CODEWRD_OUT_BIT_153_reg_model LDPC_DEC_CODEWRD_OUT_BIT_153;
    rand LDPC_DEC_CODEWRD_OUT_BIT_154_reg_model LDPC_DEC_CODEWRD_OUT_BIT_154;
    rand LDPC_DEC_CODEWRD_OUT_BIT_155_reg_model LDPC_DEC_CODEWRD_OUT_BIT_155;
    rand LDPC_DEC_CODEWRD_OUT_BIT_156_reg_model LDPC_DEC_CODEWRD_OUT_BIT_156;
    rand LDPC_DEC_CODEWRD_OUT_BIT_157_reg_model LDPC_DEC_CODEWRD_OUT_BIT_157;
    rand LDPC_DEC_CODEWRD_OUT_BIT_158_reg_model LDPC_DEC_CODEWRD_OUT_BIT_158;
    rand LDPC_DEC_CODEWRD_OUT_BIT_159_reg_model LDPC_DEC_CODEWRD_OUT_BIT_159;
    rand LDPC_DEC_CODEWRD_OUT_BIT_160_reg_model LDPC_DEC_CODEWRD_OUT_BIT_160;
    rand LDPC_DEC_CODEWRD_OUT_BIT_161_reg_model LDPC_DEC_CODEWRD_OUT_BIT_161;
    rand LDPC_DEC_CODEWRD_OUT_BIT_162_reg_model LDPC_DEC_CODEWRD_OUT_BIT_162;
    rand LDPC_DEC_CODEWRD_OUT_BIT_163_reg_model LDPC_DEC_CODEWRD_OUT_BIT_163;
    rand LDPC_DEC_CODEWRD_OUT_BIT_164_reg_model LDPC_DEC_CODEWRD_OUT_BIT_164;
    rand LDPC_DEC_CODEWRD_OUT_BIT_165_reg_model LDPC_DEC_CODEWRD_OUT_BIT_165;
    rand LDPC_DEC_CODEWRD_OUT_BIT_166_reg_model LDPC_DEC_CODEWRD_OUT_BIT_166;
    rand LDPC_DEC_CODEWRD_OUT_BIT_167_reg_model LDPC_DEC_CODEWRD_OUT_BIT_167;
    rand LDPC_DEC_CODEWRD_OUT_BIT_168_reg_model LDPC_DEC_CODEWRD_OUT_BIT_168;
    rand LDPC_DEC_CODEWRD_OUT_BIT_169_reg_model LDPC_DEC_CODEWRD_OUT_BIT_169;
    rand LDPC_DEC_CODEWRD_OUT_BIT_170_reg_model LDPC_DEC_CODEWRD_OUT_BIT_170;
    rand LDPC_DEC_CODEWRD_OUT_BIT_171_reg_model LDPC_DEC_CODEWRD_OUT_BIT_171;
    rand LDPC_DEC_CODEWRD_OUT_BIT_172_reg_model LDPC_DEC_CODEWRD_OUT_BIT_172;
    rand LDPC_DEC_CODEWRD_OUT_BIT_173_reg_model LDPC_DEC_CODEWRD_OUT_BIT_173;
    rand LDPC_DEC_CODEWRD_OUT_BIT_174_reg_model LDPC_DEC_CODEWRD_OUT_BIT_174;
    rand LDPC_DEC_CODEWRD_OUT_BIT_175_reg_model LDPC_DEC_CODEWRD_OUT_BIT_175;
    rand LDPC_DEC_CODEWRD_OUT_BIT_176_reg_model LDPC_DEC_CODEWRD_OUT_BIT_176;
    rand LDPC_DEC_CODEWRD_OUT_BIT_177_reg_model LDPC_DEC_CODEWRD_OUT_BIT_177;
    rand LDPC_DEC_CODEWRD_OUT_BIT_178_reg_model LDPC_DEC_CODEWRD_OUT_BIT_178;
    rand LDPC_DEC_CODEWRD_OUT_BIT_179_reg_model LDPC_DEC_CODEWRD_OUT_BIT_179;
    rand LDPC_DEC_CODEWRD_OUT_BIT_180_reg_model LDPC_DEC_CODEWRD_OUT_BIT_180;
    rand LDPC_DEC_CODEWRD_OUT_BIT_181_reg_model LDPC_DEC_CODEWRD_OUT_BIT_181;
    rand LDPC_DEC_CODEWRD_OUT_BIT_182_reg_model LDPC_DEC_CODEWRD_OUT_BIT_182;
    rand LDPC_DEC_CODEWRD_OUT_BIT_183_reg_model LDPC_DEC_CODEWRD_OUT_BIT_183;
    rand LDPC_DEC_CODEWRD_OUT_BIT_184_reg_model LDPC_DEC_CODEWRD_OUT_BIT_184;
    rand LDPC_DEC_CODEWRD_OUT_BIT_185_reg_model LDPC_DEC_CODEWRD_OUT_BIT_185;
    rand LDPC_DEC_CODEWRD_OUT_BIT_186_reg_model LDPC_DEC_CODEWRD_OUT_BIT_186;
    rand LDPC_DEC_CODEWRD_OUT_BIT_187_reg_model LDPC_DEC_CODEWRD_OUT_BIT_187;
    rand LDPC_DEC_CODEWRD_OUT_BIT_188_reg_model LDPC_DEC_CODEWRD_OUT_BIT_188;
    rand LDPC_DEC_CODEWRD_OUT_BIT_189_reg_model LDPC_DEC_CODEWRD_OUT_BIT_189;
    rand LDPC_DEC_CODEWRD_OUT_BIT_190_reg_model LDPC_DEC_CODEWRD_OUT_BIT_190;
    rand LDPC_DEC_CODEWRD_OUT_BIT_191_reg_model LDPC_DEC_CODEWRD_OUT_BIT_191;
    rand LDPC_DEC_CODEWRD_OUT_BIT_192_reg_model LDPC_DEC_CODEWRD_OUT_BIT_192;
    rand LDPC_DEC_CODEWRD_OUT_BIT_193_reg_model LDPC_DEC_CODEWRD_OUT_BIT_193;
    rand LDPC_DEC_CODEWRD_OUT_BIT_194_reg_model LDPC_DEC_CODEWRD_OUT_BIT_194;
    rand LDPC_DEC_CODEWRD_OUT_BIT_195_reg_model LDPC_DEC_CODEWRD_OUT_BIT_195;
    rand LDPC_DEC_CODEWRD_OUT_BIT_196_reg_model LDPC_DEC_CODEWRD_OUT_BIT_196;
    rand LDPC_DEC_CODEWRD_OUT_BIT_197_reg_model LDPC_DEC_CODEWRD_OUT_BIT_197;
    rand LDPC_DEC_CODEWRD_OUT_BIT_198_reg_model LDPC_DEC_CODEWRD_OUT_BIT_198;
    rand LDPC_DEC_CODEWRD_OUT_BIT_199_reg_model LDPC_DEC_CODEWRD_OUT_BIT_199;
    rand LDPC_DEC_CODEWRD_OUT_BIT_200_reg_model LDPC_DEC_CODEWRD_OUT_BIT_200;
    rand LDPC_DEC_CODEWRD_OUT_BIT_201_reg_model LDPC_DEC_CODEWRD_OUT_BIT_201;
    rand LDPC_DEC_CODEWRD_OUT_BIT_202_reg_model LDPC_DEC_CODEWRD_OUT_BIT_202;
    rand LDPC_DEC_CODEWRD_OUT_BIT_203_reg_model LDPC_DEC_CODEWRD_OUT_BIT_203;
    rand LDPC_DEC_CODEWRD_OUT_BIT_204_reg_model LDPC_DEC_CODEWRD_OUT_BIT_204;
    rand LDPC_DEC_CODEWRD_OUT_BIT_205_reg_model LDPC_DEC_CODEWRD_OUT_BIT_205;
    rand LDPC_DEC_CODEWRD_OUT_BIT_206_reg_model LDPC_DEC_CODEWRD_OUT_BIT_206;
    rand LDPC_DEC_CODEWRD_OUT_BIT_207_reg_model LDPC_DEC_CODEWRD_OUT_BIT_207;
    rand LDPC_DEC_PASS_FAIL_reg_model LDPC_DEC_PASS_FAIL;
    rand LDPC_DEC_pass_fail_decoder_reg_model LDPC_DEC_pass_fail_decoder;
    function new(string name);
      super.new(name, 4, 0);
    endfunction
    function void build();
      `rggen_ral_create_reg(LDPC_ENC_MSG_IN_0, '{}, 13'h0000, "RW", "g_LDPC_ENC_MSG_IN_0.u_register")
      `rggen_ral_create_reg(LDPC_ENC_MSG_IN_1, '{}, 13'h0004, "RW", "g_LDPC_ENC_MSG_IN_1.u_register")
      `rggen_ral_create_reg(LDPC_ENC_MSG_IN_2, '{}, 13'h0008, "RW", "g_LDPC_ENC_MSG_IN_2.u_register")
      `rggen_ral_create_reg(LDPC_ENC_MSG_IN_3, '{}, 13'h000c, "RW", "g_LDPC_ENC_MSG_IN_3.u_register")
      `rggen_ral_create_reg(LDPC_ENC_MSG_IN_4, '{}, 13'h0010, "RW", "g_LDPC_ENC_MSG_IN_4.u_register")
      `rggen_ral_create_reg(LDPC_ENC_MSG_IN_5, '{}, 13'h0014, "RW", "g_LDPC_ENC_MSG_IN_5.u_register")
      `rggen_ral_create_reg(LDPC_ENC_MSG_IN_6, '{}, 13'h0018, "RW", "g_LDPC_ENC_MSG_IN_6.u_register")
      `rggen_ral_create_reg(LDPC_ENC_MSG_IN_7, '{}, 13'h001c, "RW", "g_LDPC_ENC_MSG_IN_7.u_register")
      `rggen_ral_create_reg(LDPC_ENC_MSG_IN_8, '{}, 13'h0020, "RW", "g_LDPC_ENC_MSG_IN_8.u_register")
      `rggen_ral_create_reg(LDPC_ENC_MSG_IN_9, '{}, 13'h0024, "RW", "g_LDPC_ENC_MSG_IN_9.u_register")
      `rggen_ral_create_reg(LDPC_ENC_MSG_IN_10, '{}, 13'h0028, "RW", "g_LDPC_ENC_MSG_IN_10.u_register")
      `rggen_ral_create_reg(LDPC_ENC_MSG_IN_11, '{}, 13'h002c, "RW", "g_LDPC_ENC_MSG_IN_11.u_register")
      `rggen_ral_create_reg(LDPC_ENC_MSG_IN_12, '{}, 13'h0030, "RW", "g_LDPC_ENC_MSG_IN_12.u_register")
      `rggen_ral_create_reg(LDPC_ENC_MSG_IN_13, '{}, 13'h0034, "RW", "g_LDPC_ENC_MSG_IN_13.u_register")
      `rggen_ral_create_reg(LDPC_ENC_MSG_IN_14, '{}, 13'h0038, "RW", "g_LDPC_ENC_MSG_IN_14.u_register")
      `rggen_ral_create_reg(LDPC_ENC_MSG_IN_15, '{}, 13'h003c, "RW", "g_LDPC_ENC_MSG_IN_15.u_register")
      `rggen_ral_create_reg(LDPC_ENC_MSG_IN_16, '{}, 13'h0040, "RW", "g_LDPC_ENC_MSG_IN_16.u_register")
      `rggen_ral_create_reg(LDPC_ENC_MSG_IN_17, '{}, 13'h0044, "RW", "g_LDPC_ENC_MSG_IN_17.u_register")
      `rggen_ral_create_reg(LDPC_ENC_MSG_IN_18, '{}, 13'h0048, "RW", "g_LDPC_ENC_MSG_IN_18.u_register")
      `rggen_ral_create_reg(LDPC_ENC_MSG_IN_19, '{}, 13'h004c, "RW", "g_LDPC_ENC_MSG_IN_19.u_register")
      `rggen_ral_create_reg(LDPC_ENC_MSG_IN_20, '{}, 13'h0050, "RW", "g_LDPC_ENC_MSG_IN_20.u_register")
      `rggen_ral_create_reg(LDPC_ENC_MSG_IN_21, '{}, 13'h0054, "RW", "g_LDPC_ENC_MSG_IN_21.u_register")
      `rggen_ral_create_reg(LDPC_ENC_MSG_IN_22, '{}, 13'h0058, "RW", "g_LDPC_ENC_MSG_IN_22.u_register")
      `rggen_ral_create_reg(LDPC_ENC_MSG_IN_23, '{}, 13'h005c, "RW", "g_LDPC_ENC_MSG_IN_23.u_register")
      `rggen_ral_create_reg(LDPC_ENC_MSG_IN_24, '{}, 13'h0060, "RW", "g_LDPC_ENC_MSG_IN_24.u_register")
      `rggen_ral_create_reg(LDPC_ENC_MSG_IN_25, '{}, 13'h0064, "RW", "g_LDPC_ENC_MSG_IN_25.u_register")
      `rggen_ral_create_reg(LDPC_ENC_MSG_IN_26, '{}, 13'h0068, "RW", "g_LDPC_ENC_MSG_IN_26.u_register")
      `rggen_ral_create_reg(LDPC_ENC_MSG_IN_27, '{}, 13'h006c, "RW", "g_LDPC_ENC_MSG_IN_27.u_register")
      `rggen_ral_create_reg(LDPC_ENC_MSG_IN_28, '{}, 13'h0070, "RW", "g_LDPC_ENC_MSG_IN_28.u_register")
      `rggen_ral_create_reg(LDPC_ENC_MSG_IN_29, '{}, 13'h0074, "RW", "g_LDPC_ENC_MSG_IN_29.u_register")
      `rggen_ral_create_reg(LDPC_ENC_MSG_IN_30, '{}, 13'h0078, "RW", "g_LDPC_ENC_MSG_IN_30.u_register")
      `rggen_ral_create_reg(LDPC_ENC_MSG_IN_31, '{}, 13'h007c, "RW", "g_LDPC_ENC_MSG_IN_31.u_register")
      `rggen_ral_create_reg(LDPC_ENC_MSG_IN_32, '{}, 13'h0080, "RW", "g_LDPC_ENC_MSG_IN_32.u_register")
      `rggen_ral_create_reg(LDPC_ENC_MSG_IN_33, '{}, 13'h0084, "RW", "g_LDPC_ENC_MSG_IN_33.u_register")
      `rggen_ral_create_reg(LDPC_ENC_MSG_IN_34, '{}, 13'h0088, "RW", "g_LDPC_ENC_MSG_IN_34.u_register")
      `rggen_ral_create_reg(LDPC_ENC_MSG_IN_35, '{}, 13'h008c, "RW", "g_LDPC_ENC_MSG_IN_35.u_register")
      `rggen_ral_create_reg(LDPC_ENC_MSG_IN_36, '{}, 13'h0090, "RW", "g_LDPC_ENC_MSG_IN_36.u_register")
      `rggen_ral_create_reg(LDPC_ENC_MSG_IN_37, '{}, 13'h0094, "RW", "g_LDPC_ENC_MSG_IN_37.u_register")
      `rggen_ral_create_reg(LDPC_ENC_MSG_IN_38, '{}, 13'h0098, "RW", "g_LDPC_ENC_MSG_IN_38.u_register")
      `rggen_ral_create_reg(LDPC_ENC_MSG_IN_39, '{}, 13'h009c, "RW", "g_LDPC_ENC_MSG_IN_39.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_0, '{}, 13'h00a0, "RO", "g_LDPC_ENC_CODEWRD_OUT_0.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_1, '{}, 13'h00a4, "RO", "g_LDPC_ENC_CODEWRD_OUT_1.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_2, '{}, 13'h00a8, "RO", "g_LDPC_ENC_CODEWRD_OUT_2.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_3, '{}, 13'h00ac, "RO", "g_LDPC_ENC_CODEWRD_OUT_3.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_4, '{}, 13'h00b0, "RO", "g_LDPC_ENC_CODEWRD_OUT_4.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_5, '{}, 13'h00b4, "RO", "g_LDPC_ENC_CODEWRD_OUT_5.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_6, '{}, 13'h00b8, "RO", "g_LDPC_ENC_CODEWRD_OUT_6.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_7, '{}, 13'h00bc, "RO", "g_LDPC_ENC_CODEWRD_OUT_7.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_8, '{}, 13'h00c0, "RO", "g_LDPC_ENC_CODEWRD_OUT_8.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_9, '{}, 13'h00c4, "RO", "g_LDPC_ENC_CODEWRD_OUT_9.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_10, '{}, 13'h00c8, "RO", "g_LDPC_ENC_CODEWRD_OUT_10.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_11, '{}, 13'h00cc, "RO", "g_LDPC_ENC_CODEWRD_OUT_11.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_12, '{}, 13'h00d0, "RO", "g_LDPC_ENC_CODEWRD_OUT_12.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_13, '{}, 13'h00d4, "RO", "g_LDPC_ENC_CODEWRD_OUT_13.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_14, '{}, 13'h00d8, "RO", "g_LDPC_ENC_CODEWRD_OUT_14.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_15, '{}, 13'h00dc, "RO", "g_LDPC_ENC_CODEWRD_OUT_15.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_16, '{}, 13'h00e0, "RO", "g_LDPC_ENC_CODEWRD_OUT_16.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_17, '{}, 13'h00e4, "RO", "g_LDPC_ENC_CODEWRD_OUT_17.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_18, '{}, 13'h00e8, "RO", "g_LDPC_ENC_CODEWRD_OUT_18.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_19, '{}, 13'h00ec, "RO", "g_LDPC_ENC_CODEWRD_OUT_19.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_20, '{}, 13'h00f0, "RO", "g_LDPC_ENC_CODEWRD_OUT_20.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_21, '{}, 13'h00f4, "RO", "g_LDPC_ENC_CODEWRD_OUT_21.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_22, '{}, 13'h00f8, "RO", "g_LDPC_ENC_CODEWRD_OUT_22.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_23, '{}, 13'h00fc, "RO", "g_LDPC_ENC_CODEWRD_OUT_23.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_24, '{}, 13'h0100, "RO", "g_LDPC_ENC_CODEWRD_OUT_24.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_25, '{}, 13'h0104, "RO", "g_LDPC_ENC_CODEWRD_OUT_25.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_26, '{}, 13'h0108, "RO", "g_LDPC_ENC_CODEWRD_OUT_26.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_27, '{}, 13'h010c, "RO", "g_LDPC_ENC_CODEWRD_OUT_27.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_28, '{}, 13'h0110, "RO", "g_LDPC_ENC_CODEWRD_OUT_28.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_29, '{}, 13'h0114, "RO", "g_LDPC_ENC_CODEWRD_OUT_29.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_30, '{}, 13'h0118, "RO", "g_LDPC_ENC_CODEWRD_OUT_30.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_31, '{}, 13'h011c, "RO", "g_LDPC_ENC_CODEWRD_OUT_31.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_32, '{}, 13'h0120, "RO", "g_LDPC_ENC_CODEWRD_OUT_32.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_33, '{}, 13'h0124, "RO", "g_LDPC_ENC_CODEWRD_OUT_33.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_34, '{}, 13'h0128, "RO", "g_LDPC_ENC_CODEWRD_OUT_34.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_35, '{}, 13'h012c, "RO", "g_LDPC_ENC_CODEWRD_OUT_35.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_36, '{}, 13'h0130, "RO", "g_LDPC_ENC_CODEWRD_OUT_36.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_37, '{}, 13'h0134, "RO", "g_LDPC_ENC_CODEWRD_OUT_37.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_38, '{}, 13'h0138, "RO", "g_LDPC_ENC_CODEWRD_OUT_38.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_39, '{}, 13'h013c, "RO", "g_LDPC_ENC_CODEWRD_OUT_39.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_40, '{}, 13'h0140, "RO", "g_LDPC_ENC_CODEWRD_OUT_40.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_41, '{}, 13'h0144, "RO", "g_LDPC_ENC_CODEWRD_OUT_41.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_42, '{}, 13'h0148, "RO", "g_LDPC_ENC_CODEWRD_OUT_42.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_43, '{}, 13'h014c, "RO", "g_LDPC_ENC_CODEWRD_OUT_43.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_44, '{}, 13'h0150, "RO", "g_LDPC_ENC_CODEWRD_OUT_44.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_45, '{}, 13'h0154, "RO", "g_LDPC_ENC_CODEWRD_OUT_45.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_46, '{}, 13'h0158, "RO", "g_LDPC_ENC_CODEWRD_OUT_46.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_47, '{}, 13'h015c, "RO", "g_LDPC_ENC_CODEWRD_OUT_47.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_48, '{}, 13'h0160, "RO", "g_LDPC_ENC_CODEWRD_OUT_48.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_49, '{}, 13'h0164, "RO", "g_LDPC_ENC_CODEWRD_OUT_49.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_50, '{}, 13'h0168, "RO", "g_LDPC_ENC_CODEWRD_OUT_50.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_51, '{}, 13'h016c, "RO", "g_LDPC_ENC_CODEWRD_OUT_51.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_52, '{}, 13'h0170, "RO", "g_LDPC_ENC_CODEWRD_OUT_52.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_53, '{}, 13'h0174, "RO", "g_LDPC_ENC_CODEWRD_OUT_53.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_54, '{}, 13'h0178, "RO", "g_LDPC_ENC_CODEWRD_OUT_54.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_55, '{}, 13'h017c, "RO", "g_LDPC_ENC_CODEWRD_OUT_55.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_56, '{}, 13'h0180, "RO", "g_LDPC_ENC_CODEWRD_OUT_56.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_57, '{}, 13'h0184, "RO", "g_LDPC_ENC_CODEWRD_OUT_57.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_58, '{}, 13'h0188, "RO", "g_LDPC_ENC_CODEWRD_OUT_58.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_59, '{}, 13'h018c, "RO", "g_LDPC_ENC_CODEWRD_OUT_59.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_60, '{}, 13'h0190, "RO", "g_LDPC_ENC_CODEWRD_OUT_60.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_61, '{}, 13'h0194, "RO", "g_LDPC_ENC_CODEWRD_OUT_61.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_62, '{}, 13'h0198, "RO", "g_LDPC_ENC_CODEWRD_OUT_62.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_63, '{}, 13'h019c, "RO", "g_LDPC_ENC_CODEWRD_OUT_63.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_64, '{}, 13'h01a0, "RO", "g_LDPC_ENC_CODEWRD_OUT_64.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_65, '{}, 13'h01a4, "RO", "g_LDPC_ENC_CODEWRD_OUT_65.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_66, '{}, 13'h01a8, "RO", "g_LDPC_ENC_CODEWRD_OUT_66.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_67, '{}, 13'h01ac, "RO", "g_LDPC_ENC_CODEWRD_OUT_67.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_68, '{}, 13'h01b0, "RO", "g_LDPC_ENC_CODEWRD_OUT_68.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_69, '{}, 13'h01b4, "RO", "g_LDPC_ENC_CODEWRD_OUT_69.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_70, '{}, 13'h01b8, "RO", "g_LDPC_ENC_CODEWRD_OUT_70.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_71, '{}, 13'h01bc, "RO", "g_LDPC_ENC_CODEWRD_OUT_71.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_72, '{}, 13'h01c0, "RO", "g_LDPC_ENC_CODEWRD_OUT_72.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_73, '{}, 13'h01c4, "RO", "g_LDPC_ENC_CODEWRD_OUT_73.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_74, '{}, 13'h01c8, "RO", "g_LDPC_ENC_CODEWRD_OUT_74.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_75, '{}, 13'h01cc, "RO", "g_LDPC_ENC_CODEWRD_OUT_75.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_76, '{}, 13'h01d0, "RO", "g_LDPC_ENC_CODEWRD_OUT_76.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_77, '{}, 13'h01d4, "RO", "g_LDPC_ENC_CODEWRD_OUT_77.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_78, '{}, 13'h01d8, "RO", "g_LDPC_ENC_CODEWRD_OUT_78.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_79, '{}, 13'h01dc, "RO", "g_LDPC_ENC_CODEWRD_OUT_79.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_80, '{}, 13'h01e0, "RO", "g_LDPC_ENC_CODEWRD_OUT_80.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_81, '{}, 13'h01e4, "RO", "g_LDPC_ENC_CODEWRD_OUT_81.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_82, '{}, 13'h01e8, "RO", "g_LDPC_ENC_CODEWRD_OUT_82.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_83, '{}, 13'h01ec, "RO", "g_LDPC_ENC_CODEWRD_OUT_83.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_84, '{}, 13'h01f0, "RO", "g_LDPC_ENC_CODEWRD_OUT_84.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_85, '{}, 13'h01f4, "RO", "g_LDPC_ENC_CODEWRD_OUT_85.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_86, '{}, 13'h01f8, "RO", "g_LDPC_ENC_CODEWRD_OUT_86.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_87, '{}, 13'h01fc, "RO", "g_LDPC_ENC_CODEWRD_OUT_87.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_88, '{}, 13'h0200, "RO", "g_LDPC_ENC_CODEWRD_OUT_88.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_89, '{}, 13'h0204, "RO", "g_LDPC_ENC_CODEWRD_OUT_89.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_90, '{}, 13'h0208, "RO", "g_LDPC_ENC_CODEWRD_OUT_90.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_91, '{}, 13'h020c, "RO", "g_LDPC_ENC_CODEWRD_OUT_91.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_92, '{}, 13'h0210, "RO", "g_LDPC_ENC_CODEWRD_OUT_92.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_93, '{}, 13'h0214, "RO", "g_LDPC_ENC_CODEWRD_OUT_93.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_94, '{}, 13'h0218, "RO", "g_LDPC_ENC_CODEWRD_OUT_94.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_95, '{}, 13'h021c, "RO", "g_LDPC_ENC_CODEWRD_OUT_95.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_96, '{}, 13'h0220, "RO", "g_LDPC_ENC_CODEWRD_OUT_96.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_97, '{}, 13'h0224, "RO", "g_LDPC_ENC_CODEWRD_OUT_97.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_98, '{}, 13'h0228, "RO", "g_LDPC_ENC_CODEWRD_OUT_98.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_99, '{}, 13'h022c, "RO", "g_LDPC_ENC_CODEWRD_OUT_99.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_100, '{}, 13'h0230, "RO", "g_LDPC_ENC_CODEWRD_OUT_100.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_101, '{}, 13'h0234, "RO", "g_LDPC_ENC_CODEWRD_OUT_101.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_102, '{}, 13'h0238, "RO", "g_LDPC_ENC_CODEWRD_OUT_102.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_103, '{}, 13'h023c, "RO", "g_LDPC_ENC_CODEWRD_OUT_103.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_104, '{}, 13'h0240, "RO", "g_LDPC_ENC_CODEWRD_OUT_104.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_105, '{}, 13'h0244, "RO", "g_LDPC_ENC_CODEWRD_OUT_105.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_106, '{}, 13'h0248, "RO", "g_LDPC_ENC_CODEWRD_OUT_106.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_107, '{}, 13'h024c, "RO", "g_LDPC_ENC_CODEWRD_OUT_107.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_108, '{}, 13'h0250, "RO", "g_LDPC_ENC_CODEWRD_OUT_108.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_109, '{}, 13'h0254, "RO", "g_LDPC_ENC_CODEWRD_OUT_109.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_110, '{}, 13'h0258, "RO", "g_LDPC_ENC_CODEWRD_OUT_110.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_111, '{}, 13'h025c, "RO", "g_LDPC_ENC_CODEWRD_OUT_111.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_112, '{}, 13'h0260, "RO", "g_LDPC_ENC_CODEWRD_OUT_112.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_113, '{}, 13'h0264, "RO", "g_LDPC_ENC_CODEWRD_OUT_113.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_114, '{}, 13'h0268, "RO", "g_LDPC_ENC_CODEWRD_OUT_114.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_115, '{}, 13'h026c, "RO", "g_LDPC_ENC_CODEWRD_OUT_115.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_116, '{}, 13'h0270, "RO", "g_LDPC_ENC_CODEWRD_OUT_116.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_117, '{}, 13'h0274, "RO", "g_LDPC_ENC_CODEWRD_OUT_117.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_118, '{}, 13'h0278, "RO", "g_LDPC_ENC_CODEWRD_OUT_118.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_119, '{}, 13'h027c, "RO", "g_LDPC_ENC_CODEWRD_OUT_119.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_120, '{}, 13'h0280, "RO", "g_LDPC_ENC_CODEWRD_OUT_120.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_121, '{}, 13'h0284, "RO", "g_LDPC_ENC_CODEWRD_OUT_121.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_122, '{}, 13'h0288, "RO", "g_LDPC_ENC_CODEWRD_OUT_122.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_123, '{}, 13'h028c, "RO", "g_LDPC_ENC_CODEWRD_OUT_123.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_124, '{}, 13'h0290, "RO", "g_LDPC_ENC_CODEWRD_OUT_124.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_125, '{}, 13'h0294, "RO", "g_LDPC_ENC_CODEWRD_OUT_125.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_126, '{}, 13'h0298, "RO", "g_LDPC_ENC_CODEWRD_OUT_126.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_127, '{}, 13'h029c, "RO", "g_LDPC_ENC_CODEWRD_OUT_127.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_128, '{}, 13'h02a0, "RO", "g_LDPC_ENC_CODEWRD_OUT_128.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_129, '{}, 13'h02a4, "RO", "g_LDPC_ENC_CODEWRD_OUT_129.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_130, '{}, 13'h02a8, "RO", "g_LDPC_ENC_CODEWRD_OUT_130.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_131, '{}, 13'h02ac, "RO", "g_LDPC_ENC_CODEWRD_OUT_131.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_132, '{}, 13'h02b0, "RO", "g_LDPC_ENC_CODEWRD_OUT_132.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_133, '{}, 13'h02b4, "RO", "g_LDPC_ENC_CODEWRD_OUT_133.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_134, '{}, 13'h02b8, "RO", "g_LDPC_ENC_CODEWRD_OUT_134.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_135, '{}, 13'h02bc, "RO", "g_LDPC_ENC_CODEWRD_OUT_135.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_136, '{}, 13'h02c0, "RO", "g_LDPC_ENC_CODEWRD_OUT_136.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_137, '{}, 13'h02c4, "RO", "g_LDPC_ENC_CODEWRD_OUT_137.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_138, '{}, 13'h02c8, "RO", "g_LDPC_ENC_CODEWRD_OUT_138.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_139, '{}, 13'h02cc, "RO", "g_LDPC_ENC_CODEWRD_OUT_139.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_140, '{}, 13'h02d0, "RO", "g_LDPC_ENC_CODEWRD_OUT_140.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_141, '{}, 13'h02d4, "RO", "g_LDPC_ENC_CODEWRD_OUT_141.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_142, '{}, 13'h02d8, "RO", "g_LDPC_ENC_CODEWRD_OUT_142.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_143, '{}, 13'h02dc, "RO", "g_LDPC_ENC_CODEWRD_OUT_143.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_144, '{}, 13'h02e0, "RO", "g_LDPC_ENC_CODEWRD_OUT_144.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_145, '{}, 13'h02e4, "RO", "g_LDPC_ENC_CODEWRD_OUT_145.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_146, '{}, 13'h02e8, "RO", "g_LDPC_ENC_CODEWRD_OUT_146.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_147, '{}, 13'h02ec, "RO", "g_LDPC_ENC_CODEWRD_OUT_147.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_148, '{}, 13'h02f0, "RO", "g_LDPC_ENC_CODEWRD_OUT_148.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_149, '{}, 13'h02f4, "RO", "g_LDPC_ENC_CODEWRD_OUT_149.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_150, '{}, 13'h02f8, "RO", "g_LDPC_ENC_CODEWRD_OUT_150.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_151, '{}, 13'h02fc, "RO", "g_LDPC_ENC_CODEWRD_OUT_151.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_152, '{}, 13'h0300, "RO", "g_LDPC_ENC_CODEWRD_OUT_152.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_153, '{}, 13'h0304, "RO", "g_LDPC_ENC_CODEWRD_OUT_153.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_154, '{}, 13'h0308, "RO", "g_LDPC_ENC_CODEWRD_OUT_154.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_155, '{}, 13'h030c, "RO", "g_LDPC_ENC_CODEWRD_OUT_155.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_156, '{}, 13'h0310, "RO", "g_LDPC_ENC_CODEWRD_OUT_156.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_157, '{}, 13'h0314, "RO", "g_LDPC_ENC_CODEWRD_OUT_157.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_158, '{}, 13'h0318, "RO", "g_LDPC_ENC_CODEWRD_OUT_158.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_159, '{}, 13'h031c, "RO", "g_LDPC_ENC_CODEWRD_OUT_159.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_160, '{}, 13'h0320, "RO", "g_LDPC_ENC_CODEWRD_OUT_160.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_161, '{}, 13'h0324, "RO", "g_LDPC_ENC_CODEWRD_OUT_161.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_162, '{}, 13'h0328, "RO", "g_LDPC_ENC_CODEWRD_OUT_162.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_163, '{}, 13'h032c, "RO", "g_LDPC_ENC_CODEWRD_OUT_163.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_164, '{}, 13'h0330, "RO", "g_LDPC_ENC_CODEWRD_OUT_164.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_165, '{}, 13'h0334, "RO", "g_LDPC_ENC_CODEWRD_OUT_165.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_166, '{}, 13'h0338, "RO", "g_LDPC_ENC_CODEWRD_OUT_166.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_167, '{}, 13'h033c, "RO", "g_LDPC_ENC_CODEWRD_OUT_167.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_168, '{}, 13'h0340, "RO", "g_LDPC_ENC_CODEWRD_OUT_168.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_169, '{}, 13'h0344, "RO", "g_LDPC_ENC_CODEWRD_OUT_169.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_170, '{}, 13'h0348, "RO", "g_LDPC_ENC_CODEWRD_OUT_170.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_171, '{}, 13'h034c, "RO", "g_LDPC_ENC_CODEWRD_OUT_171.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_172, '{}, 13'h0350, "RO", "g_LDPC_ENC_CODEWRD_OUT_172.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_173, '{}, 13'h0354, "RO", "g_LDPC_ENC_CODEWRD_OUT_173.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_174, '{}, 13'h0358, "RO", "g_LDPC_ENC_CODEWRD_OUT_174.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_175, '{}, 13'h035c, "RO", "g_LDPC_ENC_CODEWRD_OUT_175.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_176, '{}, 13'h0360, "RO", "g_LDPC_ENC_CODEWRD_OUT_176.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_177, '{}, 13'h0364, "RO", "g_LDPC_ENC_CODEWRD_OUT_177.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_178, '{}, 13'h0368, "RO", "g_LDPC_ENC_CODEWRD_OUT_178.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_179, '{}, 13'h036c, "RO", "g_LDPC_ENC_CODEWRD_OUT_179.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_180, '{}, 13'h0370, "RO", "g_LDPC_ENC_CODEWRD_OUT_180.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_181, '{}, 13'h0374, "RO", "g_LDPC_ENC_CODEWRD_OUT_181.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_182, '{}, 13'h0378, "RO", "g_LDPC_ENC_CODEWRD_OUT_182.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_183, '{}, 13'h037c, "RO", "g_LDPC_ENC_CODEWRD_OUT_183.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_184, '{}, 13'h0380, "RO", "g_LDPC_ENC_CODEWRD_OUT_184.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_185, '{}, 13'h0384, "RO", "g_LDPC_ENC_CODEWRD_OUT_185.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_186, '{}, 13'h0388, "RO", "g_LDPC_ENC_CODEWRD_OUT_186.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_187, '{}, 13'h038c, "RO", "g_LDPC_ENC_CODEWRD_OUT_187.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_188, '{}, 13'h0390, "RO", "g_LDPC_ENC_CODEWRD_OUT_188.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_189, '{}, 13'h0394, "RO", "g_LDPC_ENC_CODEWRD_OUT_189.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_190, '{}, 13'h0398, "RO", "g_LDPC_ENC_CODEWRD_OUT_190.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_191, '{}, 13'h039c, "RO", "g_LDPC_ENC_CODEWRD_OUT_191.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_192, '{}, 13'h03a0, "RO", "g_LDPC_ENC_CODEWRD_OUT_192.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_193, '{}, 13'h03a4, "RO", "g_LDPC_ENC_CODEWRD_OUT_193.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_194, '{}, 13'h03a8, "RO", "g_LDPC_ENC_CODEWRD_OUT_194.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_195, '{}, 13'h03ac, "RO", "g_LDPC_ENC_CODEWRD_OUT_195.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_196, '{}, 13'h03b0, "RO", "g_LDPC_ENC_CODEWRD_OUT_196.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_197, '{}, 13'h03b4, "RO", "g_LDPC_ENC_CODEWRD_OUT_197.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_198, '{}, 13'h03b8, "RO", "g_LDPC_ENC_CODEWRD_OUT_198.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_199, '{}, 13'h03bc, "RO", "g_LDPC_ENC_CODEWRD_OUT_199.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_200, '{}, 13'h03c0, "RO", "g_LDPC_ENC_CODEWRD_OUT_200.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_201, '{}, 13'h03c4, "RO", "g_LDPC_ENC_CODEWRD_OUT_201.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_202, '{}, 13'h03c8, "RO", "g_LDPC_ENC_CODEWRD_OUT_202.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_203, '{}, 13'h03cc, "RO", "g_LDPC_ENC_CODEWRD_OUT_203.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_204, '{}, 13'h03d0, "RO", "g_LDPC_ENC_CODEWRD_OUT_204.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_205, '{}, 13'h03d4, "RO", "g_LDPC_ENC_CODEWRD_OUT_205.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_206, '{}, 13'h03d8, "RO", "g_LDPC_ENC_CODEWRD_OUT_206.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_OUT_207, '{}, 13'h03dc, "RO", "g_LDPC_ENC_CODEWRD_OUT_207.u_register")
      `rggen_ral_create_reg(LDPC_ENC_CODEWRD_VLD, '{}, 13'h03e0, "RO", "g_LDPC_ENC_CODEWRD_VLD.u_register")
      `rggen_ral_create_reg(LDPC_DEC_SEL_FRMC, '{}, 13'h03e4, "RW", "g_LDPC_DEC_SEL_FRMC.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_0, '{}, 13'h03e8, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_0.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_1, '{}, 13'h03ec, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_1.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_2, '{}, 13'h03f0, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_2.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_3, '{}, 13'h03f4, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_3.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_4, '{}, 13'h03f8, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_4.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_5, '{}, 13'h03fc, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_5.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_6, '{}, 13'h0400, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_6.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_7, '{}, 13'h0404, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_7.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_8, '{}, 13'h0408, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_8.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_9, '{}, 13'h040c, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_9.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_10, '{}, 13'h0410, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_10.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_11, '{}, 13'h0414, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_11.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_12, '{}, 13'h0418, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_12.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_13, '{}, 13'h041c, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_13.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_14, '{}, 13'h0420, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_14.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_15, '{}, 13'h0424, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_15.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_16, '{}, 13'h0428, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_16.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_17, '{}, 13'h042c, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_17.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_18, '{}, 13'h0430, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_18.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_19, '{}, 13'h0434, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_19.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_20, '{}, 13'h0438, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_20.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_21, '{}, 13'h043c, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_21.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_22, '{}, 13'h0440, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_22.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_23, '{}, 13'h0444, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_23.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_24, '{}, 13'h0448, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_24.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_25, '{}, 13'h044c, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_25.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_26, '{}, 13'h0450, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_26.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_27, '{}, 13'h0454, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_27.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_28, '{}, 13'h0458, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_28.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_29, '{}, 13'h045c, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_29.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_30, '{}, 13'h0460, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_30.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_31, '{}, 13'h0464, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_31.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_32, '{}, 13'h0468, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_32.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_33, '{}, 13'h046c, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_33.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_34, '{}, 13'h0470, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_34.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_35, '{}, 13'h0474, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_35.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_36, '{}, 13'h0478, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_36.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_37, '{}, 13'h047c, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_37.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_38, '{}, 13'h0480, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_38.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_39, '{}, 13'h0484, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_39.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_40, '{}, 13'h0488, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_40.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_41, '{}, 13'h048c, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_41.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_42, '{}, 13'h0490, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_42.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_43, '{}, 13'h0494, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_43.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_44, '{}, 13'h0498, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_44.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_45, '{}, 13'h049c, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_45.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_46, '{}, 13'h04a0, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_46.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_47, '{}, 13'h04a4, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_47.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_48, '{}, 13'h04a8, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_48.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_49, '{}, 13'h04ac, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_49.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_50, '{}, 13'h04b0, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_50.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_51, '{}, 13'h04b4, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_51.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_52, '{}, 13'h04b8, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_52.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_53, '{}, 13'h04bc, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_53.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_54, '{}, 13'h04c0, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_54.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_55, '{}, 13'h04c4, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_55.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_56, '{}, 13'h04c8, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_56.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_57, '{}, 13'h04cc, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_57.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_58, '{}, 13'h04d0, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_58.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_59, '{}, 13'h04d4, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_59.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_60, '{}, 13'h04d8, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_60.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_61, '{}, 13'h04dc, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_61.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_62, '{}, 13'h04e0, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_62.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_63, '{}, 13'h04e4, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_63.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_64, '{}, 13'h04e8, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_64.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_65, '{}, 13'h04ec, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_65.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_66, '{}, 13'h04f0, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_66.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_67, '{}, 13'h04f4, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_67.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_68, '{}, 13'h04f8, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_68.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_69, '{}, 13'h04fc, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_69.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_70, '{}, 13'h0500, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_70.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_71, '{}, 13'h0504, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_71.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_72, '{}, 13'h0508, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_72.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_73, '{}, 13'h050c, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_73.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_74, '{}, 13'h0510, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_74.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_75, '{}, 13'h0514, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_75.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_76, '{}, 13'h0518, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_76.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_77, '{}, 13'h051c, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_77.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_78, '{}, 13'h0520, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_78.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_79, '{}, 13'h0524, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_79.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_80, '{}, 13'h0528, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_80.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_81, '{}, 13'h052c, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_81.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_82, '{}, 13'h0530, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_82.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_83, '{}, 13'h0534, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_83.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_84, '{}, 13'h0538, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_84.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_85, '{}, 13'h053c, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_85.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_86, '{}, 13'h0540, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_86.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_87, '{}, 13'h0544, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_87.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_88, '{}, 13'h0548, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_88.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_89, '{}, 13'h054c, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_89.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_90, '{}, 13'h0550, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_90.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_91, '{}, 13'h0554, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_91.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_92, '{}, 13'h0558, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_92.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_93, '{}, 13'h055c, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_93.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_94, '{}, 13'h0560, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_94.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_95, '{}, 13'h0564, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_95.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_96, '{}, 13'h0568, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_96.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_97, '{}, 13'h056c, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_97.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_98, '{}, 13'h0570, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_98.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_99, '{}, 13'h0574, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_99.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_100, '{}, 13'h0578, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_100.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_101, '{}, 13'h057c, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_101.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_102, '{}, 13'h0580, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_102.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_103, '{}, 13'h0584, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_103.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_104, '{}, 13'h0588, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_104.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_105, '{}, 13'h058c, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_105.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_106, '{}, 13'h0590, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_106.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_107, '{}, 13'h0594, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_107.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_108, '{}, 13'h0598, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_108.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_109, '{}, 13'h059c, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_109.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_110, '{}, 13'h05a0, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_110.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_111, '{}, 13'h05a4, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_111.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_112, '{}, 13'h05a8, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_112.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_113, '{}, 13'h05ac, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_113.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_114, '{}, 13'h05b0, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_114.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_115, '{}, 13'h05b4, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_115.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_116, '{}, 13'h05b8, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_116.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_117, '{}, 13'h05bc, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_117.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_118, '{}, 13'h05c0, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_118.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_119, '{}, 13'h05c4, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_119.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_120, '{}, 13'h05c8, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_120.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_121, '{}, 13'h05cc, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_121.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_122, '{}, 13'h05d0, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_122.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_123, '{}, 13'h05d4, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_123.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_124, '{}, 13'h05d8, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_124.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_125, '{}, 13'h05dc, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_125.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_126, '{}, 13'h05e0, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_126.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_127, '{}, 13'h05e4, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_127.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_128, '{}, 13'h05e8, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_128.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_129, '{}, 13'h05ec, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_129.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_130, '{}, 13'h05f0, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_130.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_131, '{}, 13'h05f4, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_131.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_132, '{}, 13'h05f8, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_132.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_133, '{}, 13'h05fc, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_133.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_134, '{}, 13'h0600, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_134.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_135, '{}, 13'h0604, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_135.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_136, '{}, 13'h0608, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_136.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_137, '{}, 13'h060c, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_137.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_138, '{}, 13'h0610, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_138.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_139, '{}, 13'h0614, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_139.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_140, '{}, 13'h0618, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_140.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_141, '{}, 13'h061c, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_141.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_142, '{}, 13'h0620, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_142.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_143, '{}, 13'h0624, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_143.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_144, '{}, 13'h0628, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_144.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_145, '{}, 13'h062c, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_145.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_146, '{}, 13'h0630, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_146.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_147, '{}, 13'h0634, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_147.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_148, '{}, 13'h0638, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_148.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_149, '{}, 13'h063c, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_149.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_150, '{}, 13'h0640, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_150.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_151, '{}, 13'h0644, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_151.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_152, '{}, 13'h0648, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_152.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_153, '{}, 13'h064c, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_153.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_154, '{}, 13'h0650, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_154.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_155, '{}, 13'h0654, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_155.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_156, '{}, 13'h0658, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_156.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_157, '{}, 13'h065c, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_157.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_158, '{}, 13'h0660, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_158.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_159, '{}, 13'h0664, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_159.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_160, '{}, 13'h0668, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_160.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_161, '{}, 13'h066c, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_161.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_162, '{}, 13'h0670, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_162.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_163, '{}, 13'h0674, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_163.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_164, '{}, 13'h0678, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_164.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_165, '{}, 13'h067c, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_165.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_166, '{}, 13'h0680, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_166.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_167, '{}, 13'h0684, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_167.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_168, '{}, 13'h0688, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_168.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_169, '{}, 13'h068c, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_169.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_170, '{}, 13'h0690, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_170.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_171, '{}, 13'h0694, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_171.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_172, '{}, 13'h0698, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_172.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_173, '{}, 13'h069c, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_173.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_174, '{}, 13'h06a0, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_174.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_175, '{}, 13'h06a4, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_175.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_176, '{}, 13'h06a8, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_176.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_177, '{}, 13'h06ac, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_177.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_178, '{}, 13'h06b0, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_178.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_179, '{}, 13'h06b4, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_179.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_180, '{}, 13'h06b8, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_180.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_181, '{}, 13'h06bc, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_181.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_182, '{}, 13'h06c0, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_182.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_183, '{}, 13'h06c4, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_183.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_184, '{}, 13'h06c8, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_184.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_185, '{}, 13'h06cc, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_185.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_186, '{}, 13'h06d0, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_186.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_187, '{}, 13'h06d4, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_187.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_188, '{}, 13'h06d8, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_188.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_189, '{}, 13'h06dc, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_189.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_190, '{}, 13'h06e0, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_190.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_191, '{}, 13'h06e4, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_191.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_192, '{}, 13'h06e8, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_192.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_193, '{}, 13'h06ec, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_193.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_194, '{}, 13'h06f0, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_194.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_195, '{}, 13'h06f4, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_195.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_196, '{}, 13'h06f8, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_196.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_197, '{}, 13'h06fc, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_197.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_198, '{}, 13'h0700, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_198.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_199, '{}, 13'h0704, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_199.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_200, '{}, 13'h0708, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_200.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_201, '{}, 13'h070c, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_201.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_202, '{}, 13'h0710, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_202.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_203, '{}, 13'h0714, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_203.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_204, '{}, 13'h0718, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_204.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_205, '{}, 13'h071c, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_205.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_206, '{}, 13'h0720, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_206.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_0_INTRO_207, '{}, 13'h0724, "RW", "g_LDPC_DEC_ERR_Q0_0_INTRO_207.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_0, '{}, 13'h0728, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_0.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_1, '{}, 13'h072c, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_1.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_2, '{}, 13'h0730, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_2.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_3, '{}, 13'h0734, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_3.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_4, '{}, 13'h0738, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_4.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_5, '{}, 13'h073c, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_5.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_6, '{}, 13'h0740, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_6.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_7, '{}, 13'h0744, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_7.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_8, '{}, 13'h0748, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_8.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_9, '{}, 13'h074c, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_9.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_10, '{}, 13'h0750, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_10.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_11, '{}, 13'h0754, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_11.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_12, '{}, 13'h0758, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_12.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_13, '{}, 13'h075c, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_13.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_14, '{}, 13'h0760, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_14.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_15, '{}, 13'h0764, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_15.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_16, '{}, 13'h0768, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_16.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_17, '{}, 13'h076c, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_17.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_18, '{}, 13'h0770, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_18.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_19, '{}, 13'h0774, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_19.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_20, '{}, 13'h0778, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_20.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_21, '{}, 13'h077c, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_21.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_22, '{}, 13'h0780, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_22.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_23, '{}, 13'h0784, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_23.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_24, '{}, 13'h0788, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_24.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_25, '{}, 13'h078c, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_25.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_26, '{}, 13'h0790, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_26.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_27, '{}, 13'h0794, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_27.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_28, '{}, 13'h0798, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_28.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_29, '{}, 13'h079c, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_29.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_30, '{}, 13'h07a0, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_30.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_31, '{}, 13'h07a4, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_31.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_32, '{}, 13'h07a8, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_32.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_33, '{}, 13'h07ac, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_33.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_34, '{}, 13'h07b0, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_34.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_35, '{}, 13'h07b4, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_35.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_36, '{}, 13'h07b8, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_36.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_37, '{}, 13'h07bc, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_37.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_38, '{}, 13'h07c0, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_38.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_39, '{}, 13'h07c4, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_39.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_40, '{}, 13'h07c8, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_40.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_41, '{}, 13'h07cc, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_41.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_42, '{}, 13'h07d0, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_42.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_43, '{}, 13'h07d4, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_43.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_44, '{}, 13'h07d8, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_44.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_45, '{}, 13'h07dc, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_45.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_46, '{}, 13'h07e0, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_46.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_47, '{}, 13'h07e4, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_47.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_48, '{}, 13'h07e8, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_48.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_49, '{}, 13'h07ec, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_49.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_50, '{}, 13'h07f0, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_50.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_51, '{}, 13'h07f4, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_51.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_52, '{}, 13'h07f8, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_52.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_53, '{}, 13'h07fc, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_53.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_54, '{}, 13'h0800, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_54.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_55, '{}, 13'h0804, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_55.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_56, '{}, 13'h0808, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_56.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_57, '{}, 13'h080c, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_57.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_58, '{}, 13'h0810, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_58.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_59, '{}, 13'h0814, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_59.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_60, '{}, 13'h0818, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_60.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_61, '{}, 13'h081c, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_61.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_62, '{}, 13'h0820, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_62.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_63, '{}, 13'h0824, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_63.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_64, '{}, 13'h0828, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_64.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_65, '{}, 13'h082c, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_65.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_66, '{}, 13'h0830, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_66.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_67, '{}, 13'h0834, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_67.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_68, '{}, 13'h0838, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_68.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_69, '{}, 13'h083c, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_69.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_70, '{}, 13'h0840, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_70.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_71, '{}, 13'h0844, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_71.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_72, '{}, 13'h0848, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_72.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_73, '{}, 13'h084c, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_73.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_74, '{}, 13'h0850, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_74.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_75, '{}, 13'h0854, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_75.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_76, '{}, 13'h0858, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_76.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_77, '{}, 13'h085c, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_77.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_78, '{}, 13'h0860, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_78.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_79, '{}, 13'h0864, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_79.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_80, '{}, 13'h0868, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_80.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_81, '{}, 13'h086c, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_81.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_82, '{}, 13'h0870, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_82.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_83, '{}, 13'h0874, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_83.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_84, '{}, 13'h0878, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_84.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_85, '{}, 13'h087c, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_85.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_86, '{}, 13'h0880, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_86.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_87, '{}, 13'h0884, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_87.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_88, '{}, 13'h0888, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_88.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_89, '{}, 13'h088c, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_89.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_90, '{}, 13'h0890, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_90.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_91, '{}, 13'h0894, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_91.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_92, '{}, 13'h0898, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_92.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_93, '{}, 13'h089c, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_93.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_94, '{}, 13'h08a0, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_94.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_95, '{}, 13'h08a4, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_95.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_96, '{}, 13'h08a8, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_96.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_97, '{}, 13'h08ac, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_97.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_98, '{}, 13'h08b0, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_98.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_99, '{}, 13'h08b4, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_99.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_100, '{}, 13'h08b8, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_100.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_101, '{}, 13'h08bc, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_101.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_102, '{}, 13'h08c0, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_102.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_103, '{}, 13'h08c4, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_103.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_104, '{}, 13'h08c8, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_104.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_105, '{}, 13'h08cc, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_105.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_106, '{}, 13'h08d0, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_106.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_107, '{}, 13'h08d4, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_107.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_108, '{}, 13'h08d8, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_108.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_109, '{}, 13'h08dc, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_109.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_110, '{}, 13'h08e0, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_110.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_111, '{}, 13'h08e4, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_111.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_112, '{}, 13'h08e8, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_112.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_113, '{}, 13'h08ec, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_113.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_114, '{}, 13'h08f0, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_114.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_115, '{}, 13'h08f4, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_115.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_116, '{}, 13'h08f8, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_116.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_117, '{}, 13'h08fc, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_117.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_118, '{}, 13'h0900, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_118.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_119, '{}, 13'h0904, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_119.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_120, '{}, 13'h0908, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_120.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_121, '{}, 13'h090c, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_121.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_122, '{}, 13'h0910, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_122.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_123, '{}, 13'h0914, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_123.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_124, '{}, 13'h0918, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_124.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_125, '{}, 13'h091c, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_125.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_126, '{}, 13'h0920, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_126.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_127, '{}, 13'h0924, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_127.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_128, '{}, 13'h0928, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_128.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_129, '{}, 13'h092c, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_129.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_130, '{}, 13'h0930, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_130.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_131, '{}, 13'h0934, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_131.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_132, '{}, 13'h0938, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_132.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_133, '{}, 13'h093c, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_133.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_134, '{}, 13'h0940, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_134.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_135, '{}, 13'h0944, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_135.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_136, '{}, 13'h0948, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_136.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_137, '{}, 13'h094c, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_137.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_138, '{}, 13'h0950, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_138.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_139, '{}, 13'h0954, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_139.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_140, '{}, 13'h0958, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_140.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_141, '{}, 13'h095c, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_141.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_142, '{}, 13'h0960, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_142.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_143, '{}, 13'h0964, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_143.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_144, '{}, 13'h0968, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_144.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_145, '{}, 13'h096c, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_145.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_146, '{}, 13'h0970, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_146.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_147, '{}, 13'h0974, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_147.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_148, '{}, 13'h0978, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_148.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_149, '{}, 13'h097c, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_149.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_150, '{}, 13'h0980, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_150.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_151, '{}, 13'h0984, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_151.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_152, '{}, 13'h0988, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_152.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_153, '{}, 13'h098c, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_153.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_154, '{}, 13'h0990, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_154.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_155, '{}, 13'h0994, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_155.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_156, '{}, 13'h0998, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_156.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_157, '{}, 13'h099c, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_157.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_158, '{}, 13'h09a0, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_158.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_159, '{}, 13'h09a4, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_159.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_160, '{}, 13'h09a8, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_160.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_161, '{}, 13'h09ac, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_161.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_162, '{}, 13'h09b0, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_162.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_163, '{}, 13'h09b4, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_163.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_164, '{}, 13'h09b8, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_164.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_165, '{}, 13'h09bc, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_165.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_166, '{}, 13'h09c0, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_166.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_167, '{}, 13'h09c4, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_167.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_168, '{}, 13'h09c8, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_168.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_169, '{}, 13'h09cc, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_169.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_170, '{}, 13'h09d0, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_170.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_171, '{}, 13'h09d4, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_171.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_172, '{}, 13'h09d8, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_172.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_173, '{}, 13'h09dc, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_173.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_174, '{}, 13'h09e0, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_174.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_175, '{}, 13'h09e4, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_175.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_176, '{}, 13'h09e8, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_176.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_177, '{}, 13'h09ec, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_177.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_178, '{}, 13'h09f0, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_178.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_179, '{}, 13'h09f4, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_179.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_180, '{}, 13'h09f8, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_180.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_181, '{}, 13'h09fc, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_181.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_182, '{}, 13'h0a00, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_182.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_183, '{}, 13'h0a04, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_183.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_184, '{}, 13'h0a08, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_184.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_185, '{}, 13'h0a0c, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_185.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_186, '{}, 13'h0a10, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_186.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_187, '{}, 13'h0a14, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_187.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_188, '{}, 13'h0a18, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_188.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_189, '{}, 13'h0a1c, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_189.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_190, '{}, 13'h0a20, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_190.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_191, '{}, 13'h0a24, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_191.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_192, '{}, 13'h0a28, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_192.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_193, '{}, 13'h0a2c, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_193.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_194, '{}, 13'h0a30, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_194.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_195, '{}, 13'h0a34, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_195.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_196, '{}, 13'h0a38, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_196.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_197, '{}, 13'h0a3c, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_197.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_198, '{}, 13'h0a40, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_198.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_199, '{}, 13'h0a44, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_199.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_200, '{}, 13'h0a48, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_200.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_201, '{}, 13'h0a4c, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_201.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_202, '{}, 13'h0a50, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_202.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_203, '{}, 13'h0a54, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_203.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_204, '{}, 13'h0a58, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_204.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_205, '{}, 13'h0a5c, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_205.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_206, '{}, 13'h0a60, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_206.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_Q0_1_INTRO_207, '{}, 13'h0a64, "RW", "g_LDPC_DEC_ERR_Q0_1_INTRO_207.u_register")
      `rggen_ral_create_reg(LDPC_DEC_ERR_INTRODUCED, '{}, 13'h0a68, "RW", "g_LDPC_DEC_ERR_INTRODUCED.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_0, '{}, 13'h0a6c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_0.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_1, '{}, 13'h0a70, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_1.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_2, '{}, 13'h0a74, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_2.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_3, '{}, 13'h0a78, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_3.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_4, '{}, 13'h0a7c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_4.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_5, '{}, 13'h0a80, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_5.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_6, '{}, 13'h0a84, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_6.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_7, '{}, 13'h0a88, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_7.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_8, '{}, 13'h0a8c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_8.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_9, '{}, 13'h0a90, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_9.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_10, '{}, 13'h0a94, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_10.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_11, '{}, 13'h0a98, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_11.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_12, '{}, 13'h0a9c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_12.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_13, '{}, 13'h0aa0, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_13.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_14, '{}, 13'h0aa4, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_14.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_15, '{}, 13'h0aa8, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_15.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_16, '{}, 13'h0aac, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_16.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_17, '{}, 13'h0ab0, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_17.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_18, '{}, 13'h0ab4, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_18.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_19, '{}, 13'h0ab8, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_19.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_20, '{}, 13'h0abc, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_20.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_21, '{}, 13'h0ac0, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_21.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_22, '{}, 13'h0ac4, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_22.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_23, '{}, 13'h0ac8, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_23.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_24, '{}, 13'h0acc, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_24.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_25, '{}, 13'h0ad0, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_25.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_26, '{}, 13'h0ad4, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_26.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_27, '{}, 13'h0ad8, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_27.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_28, '{}, 13'h0adc, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_28.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_29, '{}, 13'h0ae0, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_29.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_30, '{}, 13'h0ae4, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_30.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_31, '{}, 13'h0ae8, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_31.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_32, '{}, 13'h0aec, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_32.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_33, '{}, 13'h0af0, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_33.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_34, '{}, 13'h0af4, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_34.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_35, '{}, 13'h0af8, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_35.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_36, '{}, 13'h0afc, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_36.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_37, '{}, 13'h0b00, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_37.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_38, '{}, 13'h0b04, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_38.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_39, '{}, 13'h0b08, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_39.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_40, '{}, 13'h0b0c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_40.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_41, '{}, 13'h0b10, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_41.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_42, '{}, 13'h0b14, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_42.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_43, '{}, 13'h0b18, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_43.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_44, '{}, 13'h0b1c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_44.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_45, '{}, 13'h0b20, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_45.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_46, '{}, 13'h0b24, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_46.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_47, '{}, 13'h0b28, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_47.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_48, '{}, 13'h0b2c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_48.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_49, '{}, 13'h0b30, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_49.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_50, '{}, 13'h0b34, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_50.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_51, '{}, 13'h0b38, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_51.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_52, '{}, 13'h0b3c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_52.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_53, '{}, 13'h0b40, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_53.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_54, '{}, 13'h0b44, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_54.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_55, '{}, 13'h0b48, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_55.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_56, '{}, 13'h0b4c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_56.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_57, '{}, 13'h0b50, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_57.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_58, '{}, 13'h0b54, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_58.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_59, '{}, 13'h0b58, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_59.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_60, '{}, 13'h0b5c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_60.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_61, '{}, 13'h0b60, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_61.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_62, '{}, 13'h0b64, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_62.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_63, '{}, 13'h0b68, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_63.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_64, '{}, 13'h0b6c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_64.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_65, '{}, 13'h0b70, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_65.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_66, '{}, 13'h0b74, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_66.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_67, '{}, 13'h0b78, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_67.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_68, '{}, 13'h0b7c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_68.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_69, '{}, 13'h0b80, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_69.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_70, '{}, 13'h0b84, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_70.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_71, '{}, 13'h0b88, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_71.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_72, '{}, 13'h0b8c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_72.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_73, '{}, 13'h0b90, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_73.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_74, '{}, 13'h0b94, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_74.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_75, '{}, 13'h0b98, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_75.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_76, '{}, 13'h0b9c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_76.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_77, '{}, 13'h0ba0, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_77.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_78, '{}, 13'h0ba4, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_78.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_79, '{}, 13'h0ba8, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_79.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_80, '{}, 13'h0bac, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_80.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_81, '{}, 13'h0bb0, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_81.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_82, '{}, 13'h0bb4, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_82.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_83, '{}, 13'h0bb8, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_83.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_84, '{}, 13'h0bbc, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_84.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_85, '{}, 13'h0bc0, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_85.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_86, '{}, 13'h0bc4, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_86.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_87, '{}, 13'h0bc8, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_87.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_88, '{}, 13'h0bcc, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_88.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_89, '{}, 13'h0bd0, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_89.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_90, '{}, 13'h0bd4, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_90.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_91, '{}, 13'h0bd8, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_91.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_92, '{}, 13'h0bdc, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_92.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_93, '{}, 13'h0be0, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_93.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_94, '{}, 13'h0be4, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_94.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_95, '{}, 13'h0be8, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_95.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_96, '{}, 13'h0bec, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_96.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_97, '{}, 13'h0bf0, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_97.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_98, '{}, 13'h0bf4, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_98.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_99, '{}, 13'h0bf8, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_99.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_100, '{}, 13'h0bfc, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_100.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_101, '{}, 13'h0c00, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_101.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_102, '{}, 13'h0c04, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_102.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_103, '{}, 13'h0c08, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_103.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_104, '{}, 13'h0c0c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_104.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_105, '{}, 13'h0c10, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_105.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_106, '{}, 13'h0c14, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_106.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_107, '{}, 13'h0c18, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_107.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_108, '{}, 13'h0c1c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_108.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_109, '{}, 13'h0c20, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_109.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_110, '{}, 13'h0c24, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_110.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_111, '{}, 13'h0c28, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_111.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_112, '{}, 13'h0c2c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_112.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_113, '{}, 13'h0c30, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_113.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_114, '{}, 13'h0c34, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_114.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_115, '{}, 13'h0c38, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_115.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_116, '{}, 13'h0c3c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_116.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_117, '{}, 13'h0c40, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_117.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_118, '{}, 13'h0c44, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_118.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_119, '{}, 13'h0c48, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_119.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_120, '{}, 13'h0c4c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_120.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_121, '{}, 13'h0c50, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_121.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_122, '{}, 13'h0c54, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_122.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_123, '{}, 13'h0c58, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_123.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_124, '{}, 13'h0c5c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_124.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_125, '{}, 13'h0c60, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_125.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_126, '{}, 13'h0c64, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_126.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_127, '{}, 13'h0c68, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_127.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_128, '{}, 13'h0c6c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_128.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_129, '{}, 13'h0c70, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_129.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_130, '{}, 13'h0c74, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_130.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_131, '{}, 13'h0c78, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_131.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_132, '{}, 13'h0c7c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_132.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_133, '{}, 13'h0c80, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_133.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_134, '{}, 13'h0c84, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_134.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_135, '{}, 13'h0c88, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_135.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_136, '{}, 13'h0c8c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_136.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_137, '{}, 13'h0c90, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_137.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_138, '{}, 13'h0c94, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_138.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_139, '{}, 13'h0c98, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_139.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_140, '{}, 13'h0c9c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_140.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_141, '{}, 13'h0ca0, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_141.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_142, '{}, 13'h0ca4, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_142.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_143, '{}, 13'h0ca8, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_143.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_144, '{}, 13'h0cac, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_144.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_145, '{}, 13'h0cb0, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_145.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_146, '{}, 13'h0cb4, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_146.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_147, '{}, 13'h0cb8, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_147.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_148, '{}, 13'h0cbc, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_148.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_149, '{}, 13'h0cc0, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_149.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_150, '{}, 13'h0cc4, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_150.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_151, '{}, 13'h0cc8, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_151.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_152, '{}, 13'h0ccc, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_152.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_153, '{}, 13'h0cd0, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_153.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_154, '{}, 13'h0cd4, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_154.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_155, '{}, 13'h0cd8, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_155.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_156, '{}, 13'h0cdc, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_156.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_157, '{}, 13'h0ce0, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_157.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_158, '{}, 13'h0ce4, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_158.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_159, '{}, 13'h0ce8, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_159.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_160, '{}, 13'h0cec, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_160.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_161, '{}, 13'h0cf0, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_161.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_162, '{}, 13'h0cf4, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_162.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_163, '{}, 13'h0cf8, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_163.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_164, '{}, 13'h0cfc, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_164.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_165, '{}, 13'h0d00, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_165.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_166, '{}, 13'h0d04, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_166.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_167, '{}, 13'h0d08, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_167.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_168, '{}, 13'h0d0c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_168.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_169, '{}, 13'h0d10, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_169.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_170, '{}, 13'h0d14, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_170.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_171, '{}, 13'h0d18, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_171.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_172, '{}, 13'h0d1c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_172.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_173, '{}, 13'h0d20, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_173.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_174, '{}, 13'h0d24, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_174.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_175, '{}, 13'h0d28, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_175.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_176, '{}, 13'h0d2c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_176.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_177, '{}, 13'h0d30, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_177.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_178, '{}, 13'h0d34, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_178.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_179, '{}, 13'h0d38, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_179.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_180, '{}, 13'h0d3c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_180.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_181, '{}, 13'h0d40, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_181.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_182, '{}, 13'h0d44, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_182.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_183, '{}, 13'h0d48, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_183.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_184, '{}, 13'h0d4c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_184.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_185, '{}, 13'h0d50, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_185.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_186, '{}, 13'h0d54, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_186.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_187, '{}, 13'h0d58, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_187.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_188, '{}, 13'h0d5c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_188.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_189, '{}, 13'h0d60, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_189.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_190, '{}, 13'h0d64, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_190.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_191, '{}, 13'h0d68, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_191.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_192, '{}, 13'h0d6c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_192.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_193, '{}, 13'h0d70, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_193.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_194, '{}, 13'h0d74, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_194.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_195, '{}, 13'h0d78, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_195.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_196, '{}, 13'h0d7c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_196.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_197, '{}, 13'h0d80, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_197.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_198, '{}, 13'h0d84, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_198.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_199, '{}, 13'h0d88, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_199.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_200, '{}, 13'h0d8c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_200.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_201, '{}, 13'h0d90, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_201.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_202, '{}, 13'h0d94, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_202.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_203, '{}, 13'h0d98, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_203.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_204, '{}, 13'h0d9c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_204.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_205, '{}, 13'h0da0, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_205.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_206, '{}, 13'h0da4, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_206.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_0_207, '{}, 13'h0da8, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_0_207.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_0, '{}, 13'h0dac, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_0.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_1, '{}, 13'h0db0, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_1.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_2, '{}, 13'h0db4, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_2.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_3, '{}, 13'h0db8, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_3.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_4, '{}, 13'h0dbc, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_4.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_5, '{}, 13'h0dc0, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_5.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_6, '{}, 13'h0dc4, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_6.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_7, '{}, 13'h0dc8, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_7.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_8, '{}, 13'h0dcc, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_8.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_9, '{}, 13'h0dd0, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_9.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_10, '{}, 13'h0dd4, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_10.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_11, '{}, 13'h0dd8, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_11.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_12, '{}, 13'h0ddc, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_12.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_13, '{}, 13'h0de0, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_13.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_14, '{}, 13'h0de4, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_14.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_15, '{}, 13'h0de8, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_15.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_16, '{}, 13'h0dec, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_16.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_17, '{}, 13'h0df0, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_17.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_18, '{}, 13'h0df4, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_18.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_19, '{}, 13'h0df8, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_19.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_20, '{}, 13'h0dfc, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_20.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_21, '{}, 13'h0e00, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_21.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_22, '{}, 13'h0e04, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_22.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_23, '{}, 13'h0e08, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_23.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_24, '{}, 13'h0e0c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_24.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_25, '{}, 13'h0e10, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_25.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_26, '{}, 13'h0e14, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_26.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_27, '{}, 13'h0e18, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_27.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_28, '{}, 13'h0e1c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_28.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_29, '{}, 13'h0e20, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_29.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_30, '{}, 13'h0e24, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_30.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_31, '{}, 13'h0e28, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_31.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_32, '{}, 13'h0e2c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_32.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_33, '{}, 13'h0e30, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_33.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_34, '{}, 13'h0e34, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_34.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_35, '{}, 13'h0e38, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_35.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_36, '{}, 13'h0e3c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_36.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_37, '{}, 13'h0e40, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_37.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_38, '{}, 13'h0e44, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_38.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_39, '{}, 13'h0e48, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_39.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_40, '{}, 13'h0e4c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_40.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_41, '{}, 13'h0e50, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_41.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_42, '{}, 13'h0e54, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_42.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_43, '{}, 13'h0e58, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_43.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_44, '{}, 13'h0e5c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_44.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_45, '{}, 13'h0e60, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_45.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_46, '{}, 13'h0e64, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_46.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_47, '{}, 13'h0e68, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_47.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_48, '{}, 13'h0e6c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_48.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_49, '{}, 13'h0e70, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_49.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_50, '{}, 13'h0e74, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_50.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_51, '{}, 13'h0e78, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_51.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_52, '{}, 13'h0e7c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_52.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_53, '{}, 13'h0e80, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_53.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_54, '{}, 13'h0e84, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_54.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_55, '{}, 13'h0e88, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_55.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_56, '{}, 13'h0e8c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_56.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_57, '{}, 13'h0e90, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_57.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_58, '{}, 13'h0e94, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_58.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_59, '{}, 13'h0e98, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_59.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_60, '{}, 13'h0e9c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_60.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_61, '{}, 13'h0ea0, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_61.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_62, '{}, 13'h0ea4, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_62.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_63, '{}, 13'h0ea8, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_63.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_64, '{}, 13'h0eac, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_64.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_65, '{}, 13'h0eb0, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_65.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_66, '{}, 13'h0eb4, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_66.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_67, '{}, 13'h0eb8, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_67.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_68, '{}, 13'h0ebc, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_68.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_69, '{}, 13'h0ec0, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_69.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_70, '{}, 13'h0ec4, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_70.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_71, '{}, 13'h0ec8, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_71.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_72, '{}, 13'h0ecc, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_72.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_73, '{}, 13'h0ed0, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_73.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_74, '{}, 13'h0ed4, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_74.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_75, '{}, 13'h0ed8, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_75.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_76, '{}, 13'h0edc, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_76.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_77, '{}, 13'h0ee0, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_77.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_78, '{}, 13'h0ee4, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_78.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_79, '{}, 13'h0ee8, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_79.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_80, '{}, 13'h0eec, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_80.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_81, '{}, 13'h0ef0, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_81.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_82, '{}, 13'h0ef4, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_82.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_83, '{}, 13'h0ef8, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_83.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_84, '{}, 13'h0efc, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_84.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_85, '{}, 13'h0f00, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_85.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_86, '{}, 13'h0f04, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_86.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_87, '{}, 13'h0f08, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_87.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_88, '{}, 13'h0f0c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_88.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_89, '{}, 13'h0f10, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_89.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_90, '{}, 13'h0f14, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_90.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_91, '{}, 13'h0f18, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_91.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_92, '{}, 13'h0f1c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_92.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_93, '{}, 13'h0f20, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_93.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_94, '{}, 13'h0f24, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_94.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_95, '{}, 13'h0f28, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_95.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_96, '{}, 13'h0f2c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_96.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_97, '{}, 13'h0f30, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_97.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_98, '{}, 13'h0f34, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_98.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_99, '{}, 13'h0f38, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_99.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_100, '{}, 13'h0f3c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_100.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_101, '{}, 13'h0f40, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_101.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_102, '{}, 13'h0f44, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_102.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_103, '{}, 13'h0f48, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_103.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_104, '{}, 13'h0f4c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_104.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_105, '{}, 13'h0f50, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_105.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_106, '{}, 13'h0f54, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_106.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_107, '{}, 13'h0f58, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_107.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_108, '{}, 13'h0f5c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_108.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_109, '{}, 13'h0f60, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_109.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_110, '{}, 13'h0f64, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_110.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_111, '{}, 13'h0f68, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_111.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_112, '{}, 13'h0f6c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_112.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_113, '{}, 13'h0f70, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_113.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_114, '{}, 13'h0f74, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_114.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_115, '{}, 13'h0f78, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_115.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_116, '{}, 13'h0f7c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_116.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_117, '{}, 13'h0f80, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_117.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_118, '{}, 13'h0f84, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_118.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_119, '{}, 13'h0f88, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_119.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_120, '{}, 13'h0f8c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_120.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_121, '{}, 13'h0f90, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_121.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_122, '{}, 13'h0f94, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_122.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_123, '{}, 13'h0f98, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_123.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_124, '{}, 13'h0f9c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_124.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_125, '{}, 13'h0fa0, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_125.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_126, '{}, 13'h0fa4, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_126.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_127, '{}, 13'h0fa8, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_127.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_128, '{}, 13'h0fac, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_128.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_129, '{}, 13'h0fb0, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_129.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_130, '{}, 13'h0fb4, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_130.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_131, '{}, 13'h0fb8, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_131.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_132, '{}, 13'h0fbc, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_132.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_133, '{}, 13'h0fc0, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_133.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_134, '{}, 13'h0fc4, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_134.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_135, '{}, 13'h0fc8, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_135.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_136, '{}, 13'h0fcc, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_136.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_137, '{}, 13'h0fd0, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_137.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_138, '{}, 13'h0fd4, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_138.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_139, '{}, 13'h0fd8, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_139.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_140, '{}, 13'h0fdc, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_140.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_141, '{}, 13'h0fe0, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_141.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_142, '{}, 13'h0fe4, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_142.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_143, '{}, 13'h0fe8, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_143.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_144, '{}, 13'h0fec, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_144.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_145, '{}, 13'h0ff0, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_145.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_146, '{}, 13'h0ff4, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_146.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_147, '{}, 13'h0ff8, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_147.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_148, '{}, 13'h0ffc, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_148.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_149, '{}, 13'h1000, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_149.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_150, '{}, 13'h1004, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_150.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_151, '{}, 13'h1008, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_151.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_152, '{}, 13'h100c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_152.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_153, '{}, 13'h1010, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_153.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_154, '{}, 13'h1014, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_154.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_155, '{}, 13'h1018, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_155.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_156, '{}, 13'h101c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_156.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_157, '{}, 13'h1020, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_157.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_158, '{}, 13'h1024, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_158.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_159, '{}, 13'h1028, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_159.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_160, '{}, 13'h102c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_160.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_161, '{}, 13'h1030, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_161.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_162, '{}, 13'h1034, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_162.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_163, '{}, 13'h1038, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_163.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_164, '{}, 13'h103c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_164.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_165, '{}, 13'h1040, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_165.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_166, '{}, 13'h1044, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_166.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_167, '{}, 13'h1048, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_167.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_168, '{}, 13'h104c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_168.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_169, '{}, 13'h1050, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_169.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_170, '{}, 13'h1054, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_170.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_171, '{}, 13'h1058, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_171.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_172, '{}, 13'h105c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_172.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_173, '{}, 13'h1060, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_173.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_174, '{}, 13'h1064, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_174.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_175, '{}, 13'h1068, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_175.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_176, '{}, 13'h106c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_176.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_177, '{}, 13'h1070, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_177.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_178, '{}, 13'h1074, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_178.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_179, '{}, 13'h1078, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_179.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_180, '{}, 13'h107c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_180.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_181, '{}, 13'h1080, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_181.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_182, '{}, 13'h1084, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_182.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_183, '{}, 13'h1088, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_183.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_184, '{}, 13'h108c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_184.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_185, '{}, 13'h1090, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_185.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_186, '{}, 13'h1094, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_186.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_187, '{}, 13'h1098, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_187.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_188, '{}, 13'h109c, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_188.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_189, '{}, 13'h10a0, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_189.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_190, '{}, 13'h10a4, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_190.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_191, '{}, 13'h10a8, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_191.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_192, '{}, 13'h10ac, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_192.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_193, '{}, 13'h10b0, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_193.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_194, '{}, 13'h10b4, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_194.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_195, '{}, 13'h10b8, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_195.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_196, '{}, 13'h10bc, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_196.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_197, '{}, 13'h10c0, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_197.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_198, '{}, 13'h10c4, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_198.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_199, '{}, 13'h10c8, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_199.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_200, '{}, 13'h10cc, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_200.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_201, '{}, 13'h10d0, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_201.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_202, '{}, 13'h10d4, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_202.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_203, '{}, 13'h10d8, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_203.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_204, '{}, 13'h10dc, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_204.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_205, '{}, 13'h10e0, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_205.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_206, '{}, 13'h10e4, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_206.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_IN_q0_1_207, '{}, 13'h10e8, "RW", "g_LDPC_DEC_CODEWRD_IN_q0_1_207.u_register")
      `rggen_ral_create_reg(LDPC_DEC_err_intro_decoder, '{}, 13'h10ec, "RO", "g_LDPC_DEC_err_intro_decoder.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_0, '{}, 13'h10f0, "RW", "g_LDPC_DEC_EXPSYND_0.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_1, '{}, 13'h10f4, "RW", "g_LDPC_DEC_EXPSYND_1.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_2, '{}, 13'h10f8, "RW", "g_LDPC_DEC_EXPSYND_2.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_3, '{}, 13'h10fc, "RW", "g_LDPC_DEC_EXPSYND_3.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_4, '{}, 13'h1100, "RW", "g_LDPC_DEC_EXPSYND_4.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_5, '{}, 13'h1104, "RW", "g_LDPC_DEC_EXPSYND_5.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_6, '{}, 13'h1108, "RW", "g_LDPC_DEC_EXPSYND_6.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_7, '{}, 13'h110c, "RW", "g_LDPC_DEC_EXPSYND_7.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_8, '{}, 13'h1110, "RW", "g_LDPC_DEC_EXPSYND_8.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_9, '{}, 13'h1114, "RW", "g_LDPC_DEC_EXPSYND_9.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_10, '{}, 13'h1118, "RW", "g_LDPC_DEC_EXPSYND_10.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_11, '{}, 13'h111c, "RW", "g_LDPC_DEC_EXPSYND_11.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_12, '{}, 13'h1120, "RW", "g_LDPC_DEC_EXPSYND_12.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_13, '{}, 13'h1124, "RW", "g_LDPC_DEC_EXPSYND_13.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_14, '{}, 13'h1128, "RW", "g_LDPC_DEC_EXPSYND_14.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_15, '{}, 13'h112c, "RW", "g_LDPC_DEC_EXPSYND_15.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_16, '{}, 13'h1130, "RW", "g_LDPC_DEC_EXPSYND_16.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_17, '{}, 13'h1134, "RW", "g_LDPC_DEC_EXPSYND_17.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_18, '{}, 13'h1138, "RW", "g_LDPC_DEC_EXPSYND_18.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_19, '{}, 13'h113c, "RW", "g_LDPC_DEC_EXPSYND_19.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_20, '{}, 13'h1140, "RW", "g_LDPC_DEC_EXPSYND_20.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_21, '{}, 13'h1144, "RW", "g_LDPC_DEC_EXPSYND_21.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_22, '{}, 13'h1148, "RW", "g_LDPC_DEC_EXPSYND_22.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_23, '{}, 13'h114c, "RW", "g_LDPC_DEC_EXPSYND_23.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_24, '{}, 13'h1150, "RW", "g_LDPC_DEC_EXPSYND_24.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_25, '{}, 13'h1154, "RW", "g_LDPC_DEC_EXPSYND_25.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_26, '{}, 13'h1158, "RW", "g_LDPC_DEC_EXPSYND_26.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_27, '{}, 13'h115c, "RW", "g_LDPC_DEC_EXPSYND_27.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_28, '{}, 13'h1160, "RW", "g_LDPC_DEC_EXPSYND_28.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_29, '{}, 13'h1164, "RW", "g_LDPC_DEC_EXPSYND_29.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_30, '{}, 13'h1168, "RW", "g_LDPC_DEC_EXPSYND_30.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_31, '{}, 13'h116c, "RW", "g_LDPC_DEC_EXPSYND_31.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_32, '{}, 13'h1170, "RW", "g_LDPC_DEC_EXPSYND_32.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_33, '{}, 13'h1174, "RW", "g_LDPC_DEC_EXPSYND_33.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_34, '{}, 13'h1178, "RW", "g_LDPC_DEC_EXPSYND_34.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_35, '{}, 13'h117c, "RW", "g_LDPC_DEC_EXPSYND_35.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_36, '{}, 13'h1180, "RW", "g_LDPC_DEC_EXPSYND_36.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_37, '{}, 13'h1184, "RW", "g_LDPC_DEC_EXPSYND_37.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_38, '{}, 13'h1188, "RW", "g_LDPC_DEC_EXPSYND_38.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_39, '{}, 13'h118c, "RW", "g_LDPC_DEC_EXPSYND_39.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_40, '{}, 13'h1190, "RW", "g_LDPC_DEC_EXPSYND_40.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_41, '{}, 13'h1194, "RW", "g_LDPC_DEC_EXPSYND_41.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_42, '{}, 13'h1198, "RW", "g_LDPC_DEC_EXPSYND_42.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_43, '{}, 13'h119c, "RW", "g_LDPC_DEC_EXPSYND_43.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_44, '{}, 13'h11a0, "RW", "g_LDPC_DEC_EXPSYND_44.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_45, '{}, 13'h11a4, "RW", "g_LDPC_DEC_EXPSYND_45.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_46, '{}, 13'h11a8, "RW", "g_LDPC_DEC_EXPSYND_46.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_47, '{}, 13'h11ac, "RW", "g_LDPC_DEC_EXPSYND_47.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_48, '{}, 13'h11b0, "RW", "g_LDPC_DEC_EXPSYND_48.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_49, '{}, 13'h11b4, "RW", "g_LDPC_DEC_EXPSYND_49.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_50, '{}, 13'h11b8, "RW", "g_LDPC_DEC_EXPSYND_50.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_51, '{}, 13'h11bc, "RW", "g_LDPC_DEC_EXPSYND_51.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_52, '{}, 13'h11c0, "RW", "g_LDPC_DEC_EXPSYND_52.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_53, '{}, 13'h11c4, "RW", "g_LDPC_DEC_EXPSYND_53.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_54, '{}, 13'h11c8, "RW", "g_LDPC_DEC_EXPSYND_54.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_55, '{}, 13'h11cc, "RW", "g_LDPC_DEC_EXPSYND_55.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_56, '{}, 13'h11d0, "RW", "g_LDPC_DEC_EXPSYND_56.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_57, '{}, 13'h11d4, "RW", "g_LDPC_DEC_EXPSYND_57.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_58, '{}, 13'h11d8, "RW", "g_LDPC_DEC_EXPSYND_58.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_59, '{}, 13'h11dc, "RW", "g_LDPC_DEC_EXPSYND_59.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_60, '{}, 13'h11e0, "RW", "g_LDPC_DEC_EXPSYND_60.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_61, '{}, 13'h11e4, "RW", "g_LDPC_DEC_EXPSYND_61.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_62, '{}, 13'h11e8, "RW", "g_LDPC_DEC_EXPSYND_62.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_63, '{}, 13'h11ec, "RW", "g_LDPC_DEC_EXPSYND_63.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_64, '{}, 13'h11f0, "RW", "g_LDPC_DEC_EXPSYND_64.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_65, '{}, 13'h11f4, "RW", "g_LDPC_DEC_EXPSYND_65.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_66, '{}, 13'h11f8, "RW", "g_LDPC_DEC_EXPSYND_66.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_67, '{}, 13'h11fc, "RW", "g_LDPC_DEC_EXPSYND_67.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_68, '{}, 13'h1200, "RW", "g_LDPC_DEC_EXPSYND_68.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_69, '{}, 13'h1204, "RW", "g_LDPC_DEC_EXPSYND_69.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_70, '{}, 13'h1208, "RW", "g_LDPC_DEC_EXPSYND_70.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_71, '{}, 13'h120c, "RW", "g_LDPC_DEC_EXPSYND_71.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_72, '{}, 13'h1210, "RW", "g_LDPC_DEC_EXPSYND_72.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_73, '{}, 13'h1214, "RW", "g_LDPC_DEC_EXPSYND_73.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_74, '{}, 13'h1218, "RW", "g_LDPC_DEC_EXPSYND_74.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_75, '{}, 13'h121c, "RW", "g_LDPC_DEC_EXPSYND_75.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_76, '{}, 13'h1220, "RW", "g_LDPC_DEC_EXPSYND_76.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_77, '{}, 13'h1224, "RW", "g_LDPC_DEC_EXPSYND_77.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_78, '{}, 13'h1228, "RW", "g_LDPC_DEC_EXPSYND_78.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_79, '{}, 13'h122c, "RW", "g_LDPC_DEC_EXPSYND_79.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_80, '{}, 13'h1230, "RW", "g_LDPC_DEC_EXPSYND_80.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_81, '{}, 13'h1234, "RW", "g_LDPC_DEC_EXPSYND_81.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_82, '{}, 13'h1238, "RW", "g_LDPC_DEC_EXPSYND_82.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_83, '{}, 13'h123c, "RW", "g_LDPC_DEC_EXPSYND_83.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_84, '{}, 13'h1240, "RW", "g_LDPC_DEC_EXPSYND_84.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_85, '{}, 13'h1244, "RW", "g_LDPC_DEC_EXPSYND_85.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_86, '{}, 13'h1248, "RW", "g_LDPC_DEC_EXPSYND_86.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_87, '{}, 13'h124c, "RW", "g_LDPC_DEC_EXPSYND_87.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_88, '{}, 13'h1250, "RW", "g_LDPC_DEC_EXPSYND_88.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_89, '{}, 13'h1254, "RW", "g_LDPC_DEC_EXPSYND_89.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_90, '{}, 13'h1258, "RW", "g_LDPC_DEC_EXPSYND_90.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_91, '{}, 13'h125c, "RW", "g_LDPC_DEC_EXPSYND_91.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_92, '{}, 13'h1260, "RW", "g_LDPC_DEC_EXPSYND_92.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_93, '{}, 13'h1264, "RW", "g_LDPC_DEC_EXPSYND_93.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_94, '{}, 13'h1268, "RW", "g_LDPC_DEC_EXPSYND_94.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_95, '{}, 13'h126c, "RW", "g_LDPC_DEC_EXPSYND_95.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_96, '{}, 13'h1270, "RW", "g_LDPC_DEC_EXPSYND_96.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_97, '{}, 13'h1274, "RW", "g_LDPC_DEC_EXPSYND_97.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_98, '{}, 13'h1278, "RW", "g_LDPC_DEC_EXPSYND_98.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_99, '{}, 13'h127c, "RW", "g_LDPC_DEC_EXPSYND_99.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_100, '{}, 13'h1280, "RW", "g_LDPC_DEC_EXPSYND_100.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_101, '{}, 13'h1284, "RW", "g_LDPC_DEC_EXPSYND_101.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_102, '{}, 13'h1288, "RW", "g_LDPC_DEC_EXPSYND_102.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_103, '{}, 13'h128c, "RW", "g_LDPC_DEC_EXPSYND_103.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_104, '{}, 13'h1290, "RW", "g_LDPC_DEC_EXPSYND_104.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_105, '{}, 13'h1294, "RW", "g_LDPC_DEC_EXPSYND_105.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_106, '{}, 13'h1298, "RW", "g_LDPC_DEC_EXPSYND_106.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_107, '{}, 13'h129c, "RW", "g_LDPC_DEC_EXPSYND_107.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_108, '{}, 13'h12a0, "RW", "g_LDPC_DEC_EXPSYND_108.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_109, '{}, 13'h12a4, "RW", "g_LDPC_DEC_EXPSYND_109.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_110, '{}, 13'h12a8, "RW", "g_LDPC_DEC_EXPSYND_110.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_111, '{}, 13'h12ac, "RW", "g_LDPC_DEC_EXPSYND_111.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_112, '{}, 13'h12b0, "RW", "g_LDPC_DEC_EXPSYND_112.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_113, '{}, 13'h12b4, "RW", "g_LDPC_DEC_EXPSYND_113.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_114, '{}, 13'h12b8, "RW", "g_LDPC_DEC_EXPSYND_114.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_115, '{}, 13'h12bc, "RW", "g_LDPC_DEC_EXPSYND_115.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_116, '{}, 13'h12c0, "RW", "g_LDPC_DEC_EXPSYND_116.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_117, '{}, 13'h12c4, "RW", "g_LDPC_DEC_EXPSYND_117.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_118, '{}, 13'h12c8, "RW", "g_LDPC_DEC_EXPSYND_118.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_119, '{}, 13'h12cc, "RW", "g_LDPC_DEC_EXPSYND_119.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_120, '{}, 13'h12d0, "RW", "g_LDPC_DEC_EXPSYND_120.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_121, '{}, 13'h12d4, "RW", "g_LDPC_DEC_EXPSYND_121.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_122, '{}, 13'h12d8, "RW", "g_LDPC_DEC_EXPSYND_122.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_123, '{}, 13'h12dc, "RW", "g_LDPC_DEC_EXPSYND_123.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_124, '{}, 13'h12e0, "RW", "g_LDPC_DEC_EXPSYND_124.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_125, '{}, 13'h12e4, "RW", "g_LDPC_DEC_EXPSYND_125.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_126, '{}, 13'h12e8, "RW", "g_LDPC_DEC_EXPSYND_126.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_127, '{}, 13'h12ec, "RW", "g_LDPC_DEC_EXPSYND_127.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_128, '{}, 13'h12f0, "RW", "g_LDPC_DEC_EXPSYND_128.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_129, '{}, 13'h12f4, "RW", "g_LDPC_DEC_EXPSYND_129.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_130, '{}, 13'h12f8, "RW", "g_LDPC_DEC_EXPSYND_130.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_131, '{}, 13'h12fc, "RW", "g_LDPC_DEC_EXPSYND_131.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_132, '{}, 13'h1300, "RW", "g_LDPC_DEC_EXPSYND_132.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_133, '{}, 13'h1304, "RW", "g_LDPC_DEC_EXPSYND_133.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_134, '{}, 13'h1308, "RW", "g_LDPC_DEC_EXPSYND_134.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_135, '{}, 13'h130c, "RW", "g_LDPC_DEC_EXPSYND_135.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_136, '{}, 13'h1310, "RW", "g_LDPC_DEC_EXPSYND_136.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_137, '{}, 13'h1314, "RW", "g_LDPC_DEC_EXPSYND_137.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_138, '{}, 13'h1318, "RW", "g_LDPC_DEC_EXPSYND_138.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_139, '{}, 13'h131c, "RW", "g_LDPC_DEC_EXPSYND_139.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_140, '{}, 13'h1320, "RW", "g_LDPC_DEC_EXPSYND_140.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_141, '{}, 13'h1324, "RW", "g_LDPC_DEC_EXPSYND_141.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_142, '{}, 13'h1328, "RW", "g_LDPC_DEC_EXPSYND_142.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_143, '{}, 13'h132c, "RW", "g_LDPC_DEC_EXPSYND_143.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_144, '{}, 13'h1330, "RW", "g_LDPC_DEC_EXPSYND_144.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_145, '{}, 13'h1334, "RW", "g_LDPC_DEC_EXPSYND_145.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_146, '{}, 13'h1338, "RW", "g_LDPC_DEC_EXPSYND_146.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_147, '{}, 13'h133c, "RW", "g_LDPC_DEC_EXPSYND_147.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_148, '{}, 13'h1340, "RW", "g_LDPC_DEC_EXPSYND_148.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_149, '{}, 13'h1344, "RW", "g_LDPC_DEC_EXPSYND_149.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_150, '{}, 13'h1348, "RW", "g_LDPC_DEC_EXPSYND_150.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_151, '{}, 13'h134c, "RW", "g_LDPC_DEC_EXPSYND_151.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_152, '{}, 13'h1350, "RW", "g_LDPC_DEC_EXPSYND_152.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_153, '{}, 13'h1354, "RW", "g_LDPC_DEC_EXPSYND_153.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_154, '{}, 13'h1358, "RW", "g_LDPC_DEC_EXPSYND_154.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_155, '{}, 13'h135c, "RW", "g_LDPC_DEC_EXPSYND_155.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_156, '{}, 13'h1360, "RW", "g_LDPC_DEC_EXPSYND_156.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_157, '{}, 13'h1364, "RW", "g_LDPC_DEC_EXPSYND_157.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_158, '{}, 13'h1368, "RW", "g_LDPC_DEC_EXPSYND_158.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_159, '{}, 13'h136c, "RW", "g_LDPC_DEC_EXPSYND_159.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_160, '{}, 13'h1370, "RW", "g_LDPC_DEC_EXPSYND_160.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_161, '{}, 13'h1374, "RW", "g_LDPC_DEC_EXPSYND_161.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_162, '{}, 13'h1378, "RW", "g_LDPC_DEC_EXPSYND_162.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_163, '{}, 13'h137c, "RW", "g_LDPC_DEC_EXPSYND_163.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_164, '{}, 13'h1380, "RW", "g_LDPC_DEC_EXPSYND_164.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_165, '{}, 13'h1384, "RW", "g_LDPC_DEC_EXPSYND_165.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_166, '{}, 13'h1388, "RW", "g_LDPC_DEC_EXPSYND_166.u_register")
      `rggen_ral_create_reg(LDPC_DEC_EXPSYND_167, '{}, 13'h138c, "RW", "g_LDPC_DEC_EXPSYND_167.u_register")
      `rggen_ral_create_reg(LDPC_DEC_PROBABILITY, '{}, 13'h1390, "RW", "g_LDPC_DEC_PROBABILITY.u_register")
      `rggen_ral_create_reg(LDPC_DEC_HAMDIST_LOOP_MAX, '{}, 13'h1394, "RW", "g_LDPC_DEC_HAMDIST_LOOP_MAX.u_register")
      `rggen_ral_create_reg(LDPC_DEC_HAMDIST_LOOP_PERCENTAGE, '{}, 13'h1398, "RW", "g_LDPC_DEC_HAMDIST_LOOP_PERCENTAGE.u_register")
      `rggen_ral_create_reg(LDPC_DEC_HAMDIST_IIR1, '{}, 13'h139c, "RW", "g_LDPC_DEC_HAMDIST_IIR1.u_register")
      `rggen_ral_create_reg(LDPC_DEC_HAMDIST_IIR2_NOT_USED, '{}, 13'h13a0, "RW", "g_LDPC_DEC_HAMDIST_IIR2_NOT_USED.u_register")
      `rggen_ral_create_reg(LDPC_DEC_HAMDIST_IIR3_NOT_USED, '{}, 13'h13a4, "RW", "g_LDPC_DEC_HAMDIST_IIR3_NOT_USED.u_register")
      `rggen_ral_create_reg(LDPC_DEC_SYN_VALID_CWORD_DEC_final, '{}, 13'h13a8, "RO", "g_LDPC_DEC_SYN_VALID_CWORD_DEC_final.u_register")
      `rggen_ral_create_reg(LDPC_DEC_START_DEC, '{}, 13'h13ac, "RW", "g_LDPC_DEC_START_DEC.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CONVERGED_LOOPS_ENDED, '{}, 13'h13b0, "RO", "g_LDPC_DEC_CONVERGED_LOOPS_ENDED.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CONVERGED_PASS_FAIL, '{}, 13'h13b4, "RO", "g_LDPC_DEC_CONVERGED_PASS_FAIL.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_0, '{}, 13'h13b8, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_0.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_1, '{}, 13'h13bc, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_1.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_2, '{}, 13'h13c0, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_2.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_3, '{}, 13'h13c4, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_3.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_4, '{}, 13'h13c8, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_4.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_5, '{}, 13'h13cc, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_5.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_6, '{}, 13'h13d0, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_6.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_7, '{}, 13'h13d4, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_7.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_8, '{}, 13'h13d8, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_8.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_9, '{}, 13'h13dc, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_9.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_10, '{}, 13'h13e0, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_10.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_11, '{}, 13'h13e4, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_11.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_12, '{}, 13'h13e8, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_12.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_13, '{}, 13'h13ec, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_13.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_14, '{}, 13'h13f0, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_14.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_15, '{}, 13'h13f4, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_15.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_16, '{}, 13'h13f8, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_16.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_17, '{}, 13'h13fc, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_17.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_18, '{}, 13'h1400, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_18.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_19, '{}, 13'h1404, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_19.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_20, '{}, 13'h1408, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_20.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_21, '{}, 13'h140c, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_21.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_22, '{}, 13'h1410, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_22.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_23, '{}, 13'h1414, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_23.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_24, '{}, 13'h1418, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_24.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_25, '{}, 13'h141c, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_25.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_26, '{}, 13'h1420, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_26.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_27, '{}, 13'h1424, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_27.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_28, '{}, 13'h1428, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_28.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_29, '{}, 13'h142c, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_29.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_30, '{}, 13'h1430, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_30.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_31, '{}, 13'h1434, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_31.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_32, '{}, 13'h1438, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_32.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_33, '{}, 13'h143c, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_33.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_34, '{}, 13'h1440, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_34.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_35, '{}, 13'h1444, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_35.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_36, '{}, 13'h1448, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_36.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_37, '{}, 13'h144c, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_37.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_38, '{}, 13'h1450, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_38.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_39, '{}, 13'h1454, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_39.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_40, '{}, 13'h1458, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_40.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_41, '{}, 13'h145c, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_41.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_42, '{}, 13'h1460, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_42.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_43, '{}, 13'h1464, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_43.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_44, '{}, 13'h1468, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_44.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_45, '{}, 13'h146c, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_45.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_46, '{}, 13'h1470, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_46.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_47, '{}, 13'h1474, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_47.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_48, '{}, 13'h1478, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_48.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_49, '{}, 13'h147c, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_49.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_50, '{}, 13'h1480, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_50.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_51, '{}, 13'h1484, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_51.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_52, '{}, 13'h1488, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_52.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_53, '{}, 13'h148c, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_53.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_54, '{}, 13'h1490, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_54.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_55, '{}, 13'h1494, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_55.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_56, '{}, 13'h1498, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_56.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_57, '{}, 13'h149c, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_57.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_58, '{}, 13'h14a0, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_58.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_59, '{}, 13'h14a4, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_59.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_60, '{}, 13'h14a8, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_60.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_61, '{}, 13'h14ac, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_61.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_62, '{}, 13'h14b0, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_62.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_63, '{}, 13'h14b4, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_63.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_64, '{}, 13'h14b8, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_64.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_65, '{}, 13'h14bc, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_65.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_66, '{}, 13'h14c0, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_66.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_67, '{}, 13'h14c4, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_67.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_68, '{}, 13'h14c8, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_68.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_69, '{}, 13'h14cc, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_69.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_70, '{}, 13'h14d0, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_70.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_71, '{}, 13'h14d4, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_71.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_72, '{}, 13'h14d8, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_72.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_73, '{}, 13'h14dc, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_73.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_74, '{}, 13'h14e0, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_74.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_75, '{}, 13'h14e4, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_75.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_76, '{}, 13'h14e8, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_76.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_77, '{}, 13'h14ec, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_77.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_78, '{}, 13'h14f0, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_78.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_79, '{}, 13'h14f4, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_79.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_80, '{}, 13'h14f8, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_80.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_81, '{}, 13'h14fc, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_81.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_82, '{}, 13'h1500, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_82.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_83, '{}, 13'h1504, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_83.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_84, '{}, 13'h1508, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_84.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_85, '{}, 13'h150c, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_85.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_86, '{}, 13'h1510, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_86.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_87, '{}, 13'h1514, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_87.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_88, '{}, 13'h1518, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_88.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_89, '{}, 13'h151c, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_89.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_90, '{}, 13'h1520, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_90.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_91, '{}, 13'h1524, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_91.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_92, '{}, 13'h1528, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_92.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_93, '{}, 13'h152c, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_93.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_94, '{}, 13'h1530, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_94.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_95, '{}, 13'h1534, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_95.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_96, '{}, 13'h1538, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_96.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_97, '{}, 13'h153c, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_97.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_98, '{}, 13'h1540, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_98.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_99, '{}, 13'h1544, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_99.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_100, '{}, 13'h1548, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_100.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_101, '{}, 13'h154c, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_101.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_102, '{}, 13'h1550, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_102.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_103, '{}, 13'h1554, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_103.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_104, '{}, 13'h1558, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_104.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_105, '{}, 13'h155c, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_105.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_106, '{}, 13'h1560, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_106.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_107, '{}, 13'h1564, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_107.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_108, '{}, 13'h1568, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_108.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_109, '{}, 13'h156c, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_109.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_110, '{}, 13'h1570, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_110.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_111, '{}, 13'h1574, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_111.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_112, '{}, 13'h1578, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_112.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_113, '{}, 13'h157c, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_113.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_114, '{}, 13'h1580, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_114.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_115, '{}, 13'h1584, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_115.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_116, '{}, 13'h1588, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_116.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_117, '{}, 13'h158c, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_117.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_118, '{}, 13'h1590, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_118.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_119, '{}, 13'h1594, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_119.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_120, '{}, 13'h1598, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_120.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_121, '{}, 13'h159c, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_121.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_122, '{}, 13'h15a0, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_122.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_123, '{}, 13'h15a4, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_123.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_124, '{}, 13'h15a8, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_124.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_125, '{}, 13'h15ac, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_125.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_126, '{}, 13'h15b0, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_126.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_127, '{}, 13'h15b4, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_127.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_128, '{}, 13'h15b8, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_128.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_129, '{}, 13'h15bc, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_129.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_130, '{}, 13'h15c0, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_130.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_131, '{}, 13'h15c4, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_131.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_132, '{}, 13'h15c8, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_132.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_133, '{}, 13'h15cc, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_133.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_134, '{}, 13'h15d0, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_134.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_135, '{}, 13'h15d4, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_135.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_136, '{}, 13'h15d8, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_136.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_137, '{}, 13'h15dc, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_137.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_138, '{}, 13'h15e0, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_138.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_139, '{}, 13'h15e4, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_139.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_140, '{}, 13'h15e8, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_140.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_141, '{}, 13'h15ec, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_141.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_142, '{}, 13'h15f0, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_142.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_143, '{}, 13'h15f4, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_143.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_144, '{}, 13'h15f8, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_144.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_145, '{}, 13'h15fc, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_145.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_146, '{}, 13'h1600, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_146.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_147, '{}, 13'h1604, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_147.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_148, '{}, 13'h1608, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_148.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_149, '{}, 13'h160c, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_149.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_150, '{}, 13'h1610, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_150.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_151, '{}, 13'h1614, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_151.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_152, '{}, 13'h1618, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_152.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_153, '{}, 13'h161c, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_153.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_154, '{}, 13'h1620, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_154.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_155, '{}, 13'h1624, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_155.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_156, '{}, 13'h1628, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_156.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_157, '{}, 13'h162c, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_157.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_158, '{}, 13'h1630, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_158.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_159, '{}, 13'h1634, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_159.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_160, '{}, 13'h1638, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_160.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_161, '{}, 13'h163c, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_161.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_162, '{}, 13'h1640, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_162.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_163, '{}, 13'h1644, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_163.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_164, '{}, 13'h1648, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_164.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_165, '{}, 13'h164c, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_165.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_166, '{}, 13'h1650, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_166.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_167, '{}, 13'h1654, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_167.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_168, '{}, 13'h1658, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_168.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_169, '{}, 13'h165c, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_169.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_170, '{}, 13'h1660, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_170.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_171, '{}, 13'h1664, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_171.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_172, '{}, 13'h1668, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_172.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_173, '{}, 13'h166c, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_173.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_174, '{}, 13'h1670, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_174.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_175, '{}, 13'h1674, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_175.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_176, '{}, 13'h1678, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_176.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_177, '{}, 13'h167c, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_177.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_178, '{}, 13'h1680, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_178.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_179, '{}, 13'h1684, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_179.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_180, '{}, 13'h1688, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_180.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_181, '{}, 13'h168c, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_181.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_182, '{}, 13'h1690, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_182.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_183, '{}, 13'h1694, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_183.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_184, '{}, 13'h1698, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_184.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_185, '{}, 13'h169c, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_185.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_186, '{}, 13'h16a0, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_186.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_187, '{}, 13'h16a4, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_187.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_188, '{}, 13'h16a8, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_188.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_189, '{}, 13'h16ac, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_189.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_190, '{}, 13'h16b0, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_190.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_191, '{}, 13'h16b4, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_191.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_192, '{}, 13'h16b8, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_192.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_193, '{}, 13'h16bc, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_193.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_194, '{}, 13'h16c0, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_194.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_195, '{}, 13'h16c4, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_195.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_196, '{}, 13'h16c8, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_196.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_197, '{}, 13'h16cc, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_197.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_198, '{}, 13'h16d0, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_198.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_199, '{}, 13'h16d4, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_199.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_200, '{}, 13'h16d8, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_200.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_201, '{}, 13'h16dc, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_201.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_202, '{}, 13'h16e0, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_202.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_203, '{}, 13'h16e4, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_203.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_204, '{}, 13'h16e8, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_204.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_205, '{}, 13'h16ec, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_205.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_206, '{}, 13'h16f0, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_206.u_register")
      `rggen_ral_create_reg(LDPC_DEC_CODEWRD_OUT_BIT_207, '{}, 13'h16f4, "RO", "g_LDPC_DEC_CODEWRD_OUT_BIT_207.u_register")
      `rggen_ral_create_reg(LDPC_DEC_PASS_FAIL, '{}, 13'h16f8, "RW", "g_LDPC_DEC_PASS_FAIL.u_register")
      `rggen_ral_create_reg(LDPC_DEC_pass_fail_decoder, '{}, 13'h16fc, "RO", "g_LDPC_DEC_pass_fail_decoder.u_register")
    endfunction
  endclass
endpackage
