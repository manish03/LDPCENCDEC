              flogtanh0x00001_0 = 
          (!flogtanh_sel[0]) ? 
                       flogtanh0x00000_0_q: 
                       flogtanh0x00000_1_q;
              flogtanh0x00001_1 = 
          (!flogtanh_sel[0]) ? 
                       flogtanh0x00000_2_q: 
                       flogtanh0x00000_3_q;
              flogtanh0x00001_2 = 
          (!flogtanh_sel[0]) ? 
                       flogtanh0x00000_4_q: 
                       flogtanh0x00000_5_q;
              flogtanh0x00001_3 = 
          (!flogtanh_sel[0]) ? 
                       flogtanh0x00000_6_q: 
                       flogtanh0x00000_7_q;
              flogtanh0x00001_4 = 
          (!flogtanh_sel[0]) ? 
                       flogtanh0x00000_8_q: 
                       flogtanh0x00000_9_q;
              flogtanh0x00001_5 = 
          (!flogtanh_sel[0]) ? 
                       flogtanh0x00000_10_q: 
                       flogtanh0x00000_11_q;
              flogtanh0x00001_6 = 
          (!flogtanh_sel[0]) ? 
                       flogtanh0x00000_12_q: 
                       flogtanh0x00000_13_q;
              flogtanh0x00001_7 = 
          (!flogtanh_sel[0]) ? 
                       flogtanh0x00000_14_q: 
                       flogtanh0x00000_15_q;
              flogtanh0x00001_8 = 
          (!flogtanh_sel[0]) ? 
                       flogtanh0x00000_16_q: 
                       flogtanh0x00000_17_q;
              flogtanh0x00001_9 = 
          (!flogtanh_sel[0]) ? 
                       flogtanh0x00000_18_q: 
                       flogtanh0x00000_19_q;
              flogtanh0x00001_10 = 
          (!flogtanh_sel[0]) ? 
                       flogtanh0x00000_20_q: 
                       flogtanh0x00000_21_q;
              flogtanh0x00001_11 = 
          (!flogtanh_sel[0]) ? 
                       flogtanh0x00000_22_q: 
                       flogtanh0x00000_23_q;
              flogtanh0x00001_12 = 
          (!flogtanh_sel[0]) ? 
                       flogtanh0x00000_24_q: 
                       flogtanh0x00000_25_q;
              flogtanh0x00001_13 = 
          (!flogtanh_sel[0]) ? 
                       flogtanh0x00000_26_q: 
                       flogtanh0x00000_27_q;
              flogtanh0x00001_14 = 
          (!flogtanh_sel[0]) ? 
                       flogtanh0x00000_28_q: 
                       flogtanh0x00000_29_q;
              flogtanh0x00001_15 = 
          (!flogtanh_sel[0]) ? 
                       flogtanh0x00000_30_q: 
                       flogtanh0x00000_31_q;
              flogtanh0x00001_16 = 
          (!flogtanh_sel[0]) ? 
                       flogtanh0x00000_32_q: 
                       flogtanh0x00000_33_q;
              flogtanh0x00001_17 = 
          (!flogtanh_sel[0]) ? 
                       flogtanh0x00000_34_q: 
                       flogtanh0x00000_35_q;
              flogtanh0x00001_18 = 
          (!flogtanh_sel[0]) ? 
                       flogtanh0x00000_36_q: 
                       flogtanh0x00000_37_q;
              flogtanh0x00001_19 = 
          (!flogtanh_sel[0]) ? 
                       flogtanh0x00000_38_q: 
                       flogtanh0x00000_39_q;
              flogtanh0x00001_20 = 
          (!flogtanh_sel[0]) ? 
                       flogtanh0x00000_40_q: 
                       flogtanh0x00000_41_q;
              flogtanh0x00001_21 = 
          (!flogtanh_sel[0]) ? 
                       flogtanh0x00000_42_q: 
                       flogtanh0x00000_43_q;
              flogtanh0x00001_22 = 
          (!flogtanh_sel[0]) ? 
                       flogtanh0x00000_44_q: 
                       flogtanh0x00000_45_q;
              flogtanh0x00001_23 = 
          (!flogtanh_sel[0]) ? 
                       flogtanh0x00000_46_q: 
                       flogtanh0x00000_47_q;
              flogtanh0x00001_24 = 
          (!flogtanh_sel[0]) ? 
                       flogtanh0x00000_48_q: 
                       flogtanh0x00000_49_q;
              flogtanh0x00001_25 = 
          (!flogtanh_sel[0]) ? 
                       flogtanh0x00000_50_q: 
                       flogtanh0x00000_51_q;
              flogtanh0x00001_26 = 
          (!flogtanh_sel[0]) ? 
                       flogtanh0x00000_52_q: 
                       flogtanh0x00000_53_q;
              flogtanh0x00001_27 = 
          (!flogtanh_sel[0]) ? 
                       flogtanh0x00000_54_q: 
                       flogtanh0x00000_55_q;
              flogtanh0x00001_28 = 
          (!flogtanh_sel[0]) ? 
                       flogtanh0x00000_56_q: 
                       flogtanh0x00000_57_q;
              flogtanh0x00001_29 = 
          (!flogtanh_sel[0]) ? 
                       flogtanh0x00000_58_q: 
                       flogtanh0x00000_59_q;
              flogtanh0x00001_30 = 
          (!flogtanh_sel[0]) ? 
                       flogtanh0x00000_60_q: 
                       flogtanh0x00000_61_q;
              flogtanh0x00001_31 = 
          (!flogtanh_sel[0]) ? 
                       flogtanh0x00000_62_q: 
                       flogtanh0x00000_63_q;
               flogtanh0x00001_32 =  flogtanh0x00000_64_q ;
              flogtanh0x00001_33 = 
          (!flogtanh_sel[0]) ? 
                       flogtanh0x00000_66_q: 
                       flogtanh0x00000_67_q;
              flogtanh0x00001_34 = 
          (!flogtanh_sel[0]) ? 
                       flogtanh0x00000_68_q: 
                       flogtanh0x00000_69_q;
              flogtanh0x00001_35 = 
          (!flogtanh_sel[0]) ? 
                       flogtanh0x00000_70_q: 
                       flogtanh0x00000_71_q;
              flogtanh0x00001_36 = 
          (!flogtanh_sel[0]) ? 
                       flogtanh0x00000_72_q: 
                       flogtanh0x00000_73_q;
              flogtanh0x00001_37 = 
          (!flogtanh_sel[0]) ? 
                       flogtanh0x00000_74_q: 
                       flogtanh0x00000_75_q;
               flogtanh0x00001_38 =  flogtanh0x00000_76_q ;
              flogtanh0x00001_39 = 
          (!flogtanh_sel[0]) ? 
                       flogtanh0x00000_78_q: 
                       flogtanh0x00000_79_q;
              flogtanh0x00001_40 = 
          (!flogtanh_sel[0]) ? 
                       flogtanh0x00000_80_q: 
                       flogtanh0x00000_81_q;
              flogtanh0x00001_41 = 
          (!flogtanh_sel[0]) ? 
                       flogtanh0x00000_82_q: 
                       flogtanh0x00000_83_q;
               flogtanh0x00001_42 =  flogtanh0x00000_84_q ;
               flogtanh0x00001_43 =  flogtanh0x00000_86_q ;
               flogtanh0x00001_44 =  flogtanh0x00000_88_q ;
               flogtanh0x00001_45 =  flogtanh0x00000_90_q ;
              flogtanh0x00001_46 = 
          (!flogtanh_sel[0]) ? 
                       flogtanh0x00000_92_q: 
                       flogtanh0x00000_93_q;
               flogtanh0x00001_47 =  flogtanh0x00000_94_q ;
               flogtanh0x00001_48 =  flogtanh0x00000_96_q ;
               flogtanh0x00001_49 =  flogtanh0x00000_98_q ;
               flogtanh0x00001_50 =  flogtanh0x00000_100_q ;
               flogtanh0x00001_51 =  flogtanh0x00000_102_q ;
              flogtanh0x00001_52 = 
          (!flogtanh_sel[0]) ? 
                       flogtanh0x00000_104_q: 
                       flogtanh0x00000_105_q;
              flogtanh0x00001_53 = 
          (!flogtanh_sel[0]) ? 
                       flogtanh0x00000_106_q: 
                       flogtanh0x00000_107_q;
               flogtanh0x00001_54 =  flogtanh0x00000_108_q ;
               flogtanh0x00001_55 =  flogtanh0x00000_110_q ;
               flogtanh0x00001_56 =  flogtanh0x00000_112_q ;
              flogtanh0x00001_57 = 
          (!flogtanh_sel[0]) ? 
                       flogtanh0x00000_114_q: 
                       flogtanh0x00000_115_q;
               flogtanh0x00001_58 =  flogtanh0x00000_116_q ;
               flogtanh0x00001_59 =  flogtanh0x00000_118_q ;
              flogtanh0x00001_60 = 
          (!flogtanh_sel[0]) ? 
                       flogtanh0x00000_120_q: 
                       flogtanh0x00000_121_q;
               flogtanh0x00001_61 =  flogtanh0x00000_122_q ;
              flogtanh0x00001_62 = 
          (!flogtanh_sel[0]) ? 
                       flogtanh0x00000_124_q: 
                       flogtanh0x00000_125_q;
               flogtanh0x00001_63 =  flogtanh0x00000_126_q ;
               flogtanh0x00001_64 =  flogtanh0x00000_128_q ;
               flogtanh0x00001_65 =  flogtanh0x00000_130_q ;
               flogtanh0x00001_66 =  flogtanh0x00000_132_q ;
               flogtanh0x00001_67 =  flogtanh0x00000_134_q ;
               flogtanh0x00001_68 =  flogtanh0x00000_136_q ;
               flogtanh0x00001_69 =  flogtanh0x00000_138_q ;
               flogtanh0x00001_70 =  flogtanh0x00000_140_q ;
               flogtanh0x00001_71 =  flogtanh0x00000_142_q ;
              flogtanh0x00001_72 = 
          (!flogtanh_sel[0]) ? 
                       flogtanh0x00000_144_q: 
                       flogtanh0x00000_145_q;
               flogtanh0x00001_73 =  flogtanh0x00000_146_q ;
               flogtanh0x00001_74 =  flogtanh0x00000_148_q ;
               flogtanh0x00001_75 =  flogtanh0x00000_150_q ;
               flogtanh0x00001_76 =  flogtanh0x00000_152_q ;
              flogtanh0x00001_77 = 
          (!flogtanh_sel[0]) ? 
                       flogtanh0x00000_154_q: 
                       flogtanh0x00000_155_q;
               flogtanh0x00001_78 =  flogtanh0x00000_156_q ;
               flogtanh0x00001_79 =  flogtanh0x00000_158_q ;
              flogtanh0x00001_80 = 
          (!flogtanh_sel[0]) ? 
                       flogtanh0x00000_160_q: 
                       flogtanh0x00000_161_q;
               flogtanh0x00001_81 =  flogtanh0x00000_162_q ;
               flogtanh0x00001_82 =  flogtanh0x00000_164_q ;
              flogtanh0x00001_83 = 
          (!flogtanh_sel[0]) ? 
                       flogtanh0x00000_166_q: 
                       flogtanh0x00000_167_q;
               flogtanh0x00001_84 =  flogtanh0x00000_168_q ;
               flogtanh0x00001_85 =  flogtanh0x00000_170_q ;
               flogtanh0x00001_86 =  flogtanh0x00000_172_q ;
               flogtanh0x00001_87 =  flogtanh0x00000_174_q ;
               flogtanh0x00001_88 =  flogtanh0x00000_176_q ;
               flogtanh0x00001_89 =  flogtanh0x00000_178_q ;
               flogtanh0x00001_90 =  flogtanh0x00000_180_q ;
               flogtanh0x00001_91 =  flogtanh0x00000_182_q ;
               flogtanh0x00001_92 =  flogtanh0x00000_184_q ;
               flogtanh0x00001_93 =  flogtanh0x00000_186_q ;
               flogtanh0x00001_94 =  flogtanh0x00000_188_q ;
              flogtanh0x00001_95 = 
          (!flogtanh_sel[0]) ? 
                       flogtanh0x00000_190_q: 
                       flogtanh0x00000_191_q;
               flogtanh0x00001_96 =  flogtanh0x00000_192_q ;
               flogtanh0x00001_97 =  flogtanh0x00000_194_q ;
               flogtanh0x00001_98 =  flogtanh0x00000_196_q ;
               flogtanh0x00001_99 =  flogtanh0x00000_198_q ;
               flogtanh0x00001_100 =  flogtanh0x00000_200_q ;
               flogtanh0x00001_101 =  flogtanh0x00000_202_q ;
               flogtanh0x00001_102 =  flogtanh0x00000_204_q ;
               flogtanh0x00001_103 =  flogtanh0x00000_206_q ;
               flogtanh0x00001_104 =  flogtanh0x00000_208_q ;
               flogtanh0x00001_105 =  flogtanh0x00000_210_q ;
               flogtanh0x00001_106 =  flogtanh0x00000_212_q ;
              flogtanh0x00001_107 = 
          (!flogtanh_sel[0]) ? 
                       flogtanh0x00000_214_q: 
                       flogtanh0x00000_215_q;
               flogtanh0x00001_108 =  flogtanh0x00000_216_q ;
               flogtanh0x00001_109 =  flogtanh0x00000_218_q ;
               flogtanh0x00001_110 =  flogtanh0x00000_220_q ;
               flogtanh0x00001_111 =  flogtanh0x00000_222_q ;
               flogtanh0x00001_112 =  flogtanh0x00000_224_q ;
               flogtanh0x00001_113 =  flogtanh0x00000_226_q ;
               flogtanh0x00001_114 =  flogtanh0x00000_228_q ;
              flogtanh0x00001_115 = 
          (!flogtanh_sel[0]) ? 
                       flogtanh0x00000_230_q: 
                       flogtanh0x00000_231_q;
               flogtanh0x00001_116 =  flogtanh0x00000_232_q ;
               flogtanh0x00001_117 =  flogtanh0x00000_234_q ;
               flogtanh0x00001_118 =  flogtanh0x00000_236_q ;
               flogtanh0x00001_119 =  flogtanh0x00000_238_q ;
               flogtanh0x00001_120 =  flogtanh0x00000_240_q ;
               flogtanh0x00001_121 =  flogtanh0x00000_242_q ;
               flogtanh0x00001_122 =  flogtanh0x00000_244_q ;
               flogtanh0x00001_123 =  flogtanh0x00000_246_q ;
               flogtanh0x00001_124 =  flogtanh0x00000_248_q ;
               flogtanh0x00001_125 =  flogtanh0x00000_250_q ;
               flogtanh0x00001_126 =  flogtanh0x00000_252_q ;
               flogtanh0x00001_127 =  flogtanh0x00000_254_q ;
               flogtanh0x00001_128 =  flogtanh0x00000_256_q ;
               flogtanh0x00001_129 =  flogtanh0x00000_258_q ;
               flogtanh0x00001_130 =  flogtanh0x00000_260_q ;
               flogtanh0x00001_131 =  flogtanh0x00000_262_q ;
               flogtanh0x00001_132 =  flogtanh0x00000_264_q ;
               flogtanh0x00001_133 =  flogtanh0x00000_266_q ;
               flogtanh0x00001_134 =  flogtanh0x00000_268_q ;
               flogtanh0x00001_135 =  flogtanh0x00000_270_q ;
               flogtanh0x00001_136 =  flogtanh0x00000_272_q ;
               flogtanh0x00001_137 =  flogtanh0x00000_274_q ;
               flogtanh0x00001_138 =  flogtanh0x00000_276_q ;
               flogtanh0x00001_139 =  flogtanh0x00000_278_q ;
               flogtanh0x00001_140 =  flogtanh0x00000_280_q ;
               flogtanh0x00001_141 =  flogtanh0x00000_282_q ;
              flogtanh0x00001_142 = 
          (!flogtanh_sel[0]) ? 
                       flogtanh0x00000_284_q: 
                       flogtanh0x00000_285_q;
               flogtanh0x00001_143 =  flogtanh0x00000_286_q ;
               flogtanh0x00001_144 =  flogtanh0x00000_288_q ;
               flogtanh0x00001_145 =  flogtanh0x00000_290_q ;
               flogtanh0x00001_146 =  flogtanh0x00000_292_q ;
               flogtanh0x00001_147 =  flogtanh0x00000_294_q ;
               flogtanh0x00001_148 =  flogtanh0x00000_296_q ;
               flogtanh0x00001_149 =  flogtanh0x00000_298_q ;
               flogtanh0x00001_150 =  flogtanh0x00000_300_q ;
               flogtanh0x00001_151 =  flogtanh0x00000_302_q ;
               flogtanh0x00001_152 =  flogtanh0x00000_304_q ;
               flogtanh0x00001_153 =  flogtanh0x00000_306_q ;
               flogtanh0x00001_154 =  flogtanh0x00000_308_q ;
               flogtanh0x00001_155 =  flogtanh0x00000_310_q ;
               flogtanh0x00001_156 =  flogtanh0x00000_312_q ;
               flogtanh0x00001_157 =  flogtanh0x00000_314_q ;
               flogtanh0x00001_158 =  flogtanh0x00000_316_q ;
               flogtanh0x00001_159 =  flogtanh0x00000_318_q ;
               flogtanh0x00001_160 =  flogtanh0x00000_320_q ;
               flogtanh0x00001_161 =  flogtanh0x00000_322_q ;
               flogtanh0x00001_162 =  flogtanh0x00000_324_q ;
               flogtanh0x00001_163 =  flogtanh0x00000_326_q ;
               flogtanh0x00001_164 =  flogtanh0x00000_328_q ;
               flogtanh0x00001_165 =  flogtanh0x00000_330_q ;
               flogtanh0x00001_166 =  flogtanh0x00000_332_q ;
               flogtanh0x00001_167 =  flogtanh0x00000_334_q ;
               flogtanh0x00001_168 =  flogtanh0x00000_336_q ;
               flogtanh0x00001_169 =  flogtanh0x00000_338_q ;
               flogtanh0x00001_170 =  flogtanh0x00000_340_q ;
               flogtanh0x00001_171 =  flogtanh0x00000_342_q ;
               flogtanh0x00001_172 =  flogtanh0x00000_344_q ;
               flogtanh0x00001_173 =  flogtanh0x00000_346_q ;
               flogtanh0x00001_174 =  flogtanh0x00000_348_q ;
               flogtanh0x00001_175 =  flogtanh0x00000_350_q ;
               flogtanh0x00001_176 =  flogtanh0x00000_352_q ;
              flogtanh0x00001_177 = 
          (!flogtanh_sel[0]) ? 
                       flogtanh0x00000_354_q: 
                       flogtanh0x00000_355_q;
