reg [flogtanh_WDTH -1:0] flogtanh0x00000_0,  flogtanh0x00000_0_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_1,  flogtanh0x00000_1_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_2,  flogtanh0x00000_2_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_3,  flogtanh0x00000_3_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_4,  flogtanh0x00000_4_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_5,  flogtanh0x00000_5_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_6,  flogtanh0x00000_6_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_7,  flogtanh0x00000_7_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_8,  flogtanh0x00000_8_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_9,  flogtanh0x00000_9_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_10,  flogtanh0x00000_10_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_11,  flogtanh0x00000_11_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_12,  flogtanh0x00000_12_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_13,  flogtanh0x00000_13_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_14,  flogtanh0x00000_14_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_15,  flogtanh0x00000_15_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_16,  flogtanh0x00000_16_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_17,  flogtanh0x00000_17_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_18,  flogtanh0x00000_18_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_19,  flogtanh0x00000_19_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_20,  flogtanh0x00000_20_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_21,  flogtanh0x00000_21_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_22,  flogtanh0x00000_22_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_23,  flogtanh0x00000_23_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_24,  flogtanh0x00000_24_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_25,  flogtanh0x00000_25_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_26,  flogtanh0x00000_26_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_27,  flogtanh0x00000_27_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_28,  flogtanh0x00000_28_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_29,  flogtanh0x00000_29_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_30,  flogtanh0x00000_30_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_31,  flogtanh0x00000_31_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_32,  flogtanh0x00000_32_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_33,  flogtanh0x00000_33_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_34,  flogtanh0x00000_34_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_35,  flogtanh0x00000_35_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_36,  flogtanh0x00000_36_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_37,  flogtanh0x00000_37_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_38,  flogtanh0x00000_38_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_39,  flogtanh0x00000_39_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_40,  flogtanh0x00000_40_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_41,  flogtanh0x00000_41_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_42,  flogtanh0x00000_42_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_43,  flogtanh0x00000_43_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_44,  flogtanh0x00000_44_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_45,  flogtanh0x00000_45_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_46,  flogtanh0x00000_46_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_47,  flogtanh0x00000_47_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_48,  flogtanh0x00000_48_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_49,  flogtanh0x00000_49_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_50,  flogtanh0x00000_50_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_51,  flogtanh0x00000_51_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_52,  flogtanh0x00000_52_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_53,  flogtanh0x00000_53_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_54,  flogtanh0x00000_54_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_55,  flogtanh0x00000_55_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_56,  flogtanh0x00000_56_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_57,  flogtanh0x00000_57_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_58,  flogtanh0x00000_58_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_59,  flogtanh0x00000_59_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_60,  flogtanh0x00000_60_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_61,  flogtanh0x00000_61_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_62,  flogtanh0x00000_62_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_63,  flogtanh0x00000_63_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_64,  flogtanh0x00000_64_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_65,  flogtanh0x00000_65_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_66,  flogtanh0x00000_66_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_67,  flogtanh0x00000_67_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_68,  flogtanh0x00000_68_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_69,  flogtanh0x00000_69_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_70,  flogtanh0x00000_70_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_71,  flogtanh0x00000_71_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_72,  flogtanh0x00000_72_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_73,  flogtanh0x00000_73_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_74,  flogtanh0x00000_74_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_75,  flogtanh0x00000_75_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_76,  flogtanh0x00000_76_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_77,  flogtanh0x00000_77_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_78,  flogtanh0x00000_78_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_79,  flogtanh0x00000_79_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_80,  flogtanh0x00000_80_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_81,  flogtanh0x00000_81_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_82,  flogtanh0x00000_82_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_83,  flogtanh0x00000_83_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_84,  flogtanh0x00000_84_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_85,  flogtanh0x00000_85_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_86,  flogtanh0x00000_86_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_87,  flogtanh0x00000_87_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_88,  flogtanh0x00000_88_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_89,  flogtanh0x00000_89_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_90,  flogtanh0x00000_90_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_91,  flogtanh0x00000_91_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_92,  flogtanh0x00000_92_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_93,  flogtanh0x00000_93_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_94,  flogtanh0x00000_94_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_95,  flogtanh0x00000_95_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_96,  flogtanh0x00000_96_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_97,  flogtanh0x00000_97_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_98,  flogtanh0x00000_98_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_99,  flogtanh0x00000_99_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_100,  flogtanh0x00000_100_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_101,  flogtanh0x00000_101_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_102,  flogtanh0x00000_102_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_103,  flogtanh0x00000_103_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_104,  flogtanh0x00000_104_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_105,  flogtanh0x00000_105_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_106,  flogtanh0x00000_106_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_107,  flogtanh0x00000_107_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_108,  flogtanh0x00000_108_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_109,  flogtanh0x00000_109_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_110,  flogtanh0x00000_110_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_111,  flogtanh0x00000_111_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_112,  flogtanh0x00000_112_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_113,  flogtanh0x00000_113_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_114,  flogtanh0x00000_114_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_115,  flogtanh0x00000_115_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_116,  flogtanh0x00000_116_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_117,  flogtanh0x00000_117_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_118,  flogtanh0x00000_118_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_119,  flogtanh0x00000_119_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_120,  flogtanh0x00000_120_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_121,  flogtanh0x00000_121_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_122,  flogtanh0x00000_122_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_123,  flogtanh0x00000_123_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_124,  flogtanh0x00000_124_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_125,  flogtanh0x00000_125_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_126,  flogtanh0x00000_126_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_127,  flogtanh0x00000_127_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_128,  flogtanh0x00000_128_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_129,  flogtanh0x00000_129_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_130,  flogtanh0x00000_130_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_131,  flogtanh0x00000_131_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_132,  flogtanh0x00000_132_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_133,  flogtanh0x00000_133_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_134,  flogtanh0x00000_134_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_135,  flogtanh0x00000_135_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_136,  flogtanh0x00000_136_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_137,  flogtanh0x00000_137_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_138,  flogtanh0x00000_138_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_139,  flogtanh0x00000_139_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_140,  flogtanh0x00000_140_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_141,  flogtanh0x00000_141_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_142,  flogtanh0x00000_142_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_143,  flogtanh0x00000_143_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_144,  flogtanh0x00000_144_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_145,  flogtanh0x00000_145_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_146,  flogtanh0x00000_146_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_147,  flogtanh0x00000_147_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_148,  flogtanh0x00000_148_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_149,  flogtanh0x00000_149_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_150,  flogtanh0x00000_150_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_151,  flogtanh0x00000_151_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_152,  flogtanh0x00000_152_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_153,  flogtanh0x00000_153_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_154,  flogtanh0x00000_154_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_155,  flogtanh0x00000_155_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_156,  flogtanh0x00000_156_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_157,  flogtanh0x00000_157_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_158,  flogtanh0x00000_158_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_159,  flogtanh0x00000_159_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_160,  flogtanh0x00000_160_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_161,  flogtanh0x00000_161_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_162,  flogtanh0x00000_162_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_163,  flogtanh0x00000_163_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_164,  flogtanh0x00000_164_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_165,  flogtanh0x00000_165_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_166,  flogtanh0x00000_166_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_167,  flogtanh0x00000_167_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_168,  flogtanh0x00000_168_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_169,  flogtanh0x00000_169_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_170,  flogtanh0x00000_170_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_171,  flogtanh0x00000_171_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_172,  flogtanh0x00000_172_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_173,  flogtanh0x00000_173_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_174,  flogtanh0x00000_174_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_175,  flogtanh0x00000_175_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_176,  flogtanh0x00000_176_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_177,  flogtanh0x00000_177_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_178,  flogtanh0x00000_178_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_179,  flogtanh0x00000_179_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_180,  flogtanh0x00000_180_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_181,  flogtanh0x00000_181_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_182,  flogtanh0x00000_182_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_183,  flogtanh0x00000_183_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_184,  flogtanh0x00000_184_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_185,  flogtanh0x00000_185_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_186,  flogtanh0x00000_186_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_187,  flogtanh0x00000_187_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_188,  flogtanh0x00000_188_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_189,  flogtanh0x00000_189_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_190,  flogtanh0x00000_190_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_191,  flogtanh0x00000_191_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_192,  flogtanh0x00000_192_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_193,  flogtanh0x00000_193_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_194,  flogtanh0x00000_194_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_195,  flogtanh0x00000_195_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_196,  flogtanh0x00000_196_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_197,  flogtanh0x00000_197_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_198,  flogtanh0x00000_198_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_199,  flogtanh0x00000_199_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_200,  flogtanh0x00000_200_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_201,  flogtanh0x00000_201_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_202,  flogtanh0x00000_202_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_203,  flogtanh0x00000_203_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_204,  flogtanh0x00000_204_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_205,  flogtanh0x00000_205_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_206,  flogtanh0x00000_206_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_207,  flogtanh0x00000_207_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_208,  flogtanh0x00000_208_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_209,  flogtanh0x00000_209_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_210,  flogtanh0x00000_210_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_211,  flogtanh0x00000_211_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_212,  flogtanh0x00000_212_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_213,  flogtanh0x00000_213_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_214,  flogtanh0x00000_214_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_215,  flogtanh0x00000_215_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_216,  flogtanh0x00000_216_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_217,  flogtanh0x00000_217_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_218,  flogtanh0x00000_218_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_219,  flogtanh0x00000_219_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_220,  flogtanh0x00000_220_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_221,  flogtanh0x00000_221_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_222,  flogtanh0x00000_222_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_223,  flogtanh0x00000_223_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_224,  flogtanh0x00000_224_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_225,  flogtanh0x00000_225_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_226,  flogtanh0x00000_226_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_227,  flogtanh0x00000_227_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_228,  flogtanh0x00000_228_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_229,  flogtanh0x00000_229_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_230,  flogtanh0x00000_230_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_231,  flogtanh0x00000_231_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_232,  flogtanh0x00000_232_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_233,  flogtanh0x00000_233_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_234,  flogtanh0x00000_234_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_235,  flogtanh0x00000_235_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_236,  flogtanh0x00000_236_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_237,  flogtanh0x00000_237_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_238,  flogtanh0x00000_238_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_239,  flogtanh0x00000_239_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_240,  flogtanh0x00000_240_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_241,  flogtanh0x00000_241_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_242,  flogtanh0x00000_242_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_243,  flogtanh0x00000_243_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_244,  flogtanh0x00000_244_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_245,  flogtanh0x00000_245_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_246,  flogtanh0x00000_246_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_247,  flogtanh0x00000_247_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_248,  flogtanh0x00000_248_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_249,  flogtanh0x00000_249_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_250,  flogtanh0x00000_250_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_251,  flogtanh0x00000_251_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_252,  flogtanh0x00000_252_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_253,  flogtanh0x00000_253_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_254,  flogtanh0x00000_254_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_255,  flogtanh0x00000_255_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_256,  flogtanh0x00000_256_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_257,  flogtanh0x00000_257_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_258,  flogtanh0x00000_258_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_259,  flogtanh0x00000_259_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_260,  flogtanh0x00000_260_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_261,  flogtanh0x00000_261_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_262,  flogtanh0x00000_262_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_263,  flogtanh0x00000_263_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_264,  flogtanh0x00000_264_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_265,  flogtanh0x00000_265_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_266,  flogtanh0x00000_266_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_267,  flogtanh0x00000_267_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_268,  flogtanh0x00000_268_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_269,  flogtanh0x00000_269_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_270,  flogtanh0x00000_270_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_271,  flogtanh0x00000_271_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_272,  flogtanh0x00000_272_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_273,  flogtanh0x00000_273_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_274,  flogtanh0x00000_274_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_275,  flogtanh0x00000_275_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_276,  flogtanh0x00000_276_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_277,  flogtanh0x00000_277_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_278,  flogtanh0x00000_278_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_279,  flogtanh0x00000_279_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_280,  flogtanh0x00000_280_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_281,  flogtanh0x00000_281_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_282,  flogtanh0x00000_282_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_283,  flogtanh0x00000_283_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_284,  flogtanh0x00000_284_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_285,  flogtanh0x00000_285_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_286,  flogtanh0x00000_286_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_287,  flogtanh0x00000_287_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_288,  flogtanh0x00000_288_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_289,  flogtanh0x00000_289_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_290,  flogtanh0x00000_290_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_291,  flogtanh0x00000_291_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_292,  flogtanh0x00000_292_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_293,  flogtanh0x00000_293_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_294,  flogtanh0x00000_294_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_295,  flogtanh0x00000_295_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_296,  flogtanh0x00000_296_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_297,  flogtanh0x00000_297_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_298,  flogtanh0x00000_298_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_299,  flogtanh0x00000_299_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_300,  flogtanh0x00000_300_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_301,  flogtanh0x00000_301_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_302,  flogtanh0x00000_302_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_303,  flogtanh0x00000_303_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_304,  flogtanh0x00000_304_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_305,  flogtanh0x00000_305_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_306,  flogtanh0x00000_306_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_307,  flogtanh0x00000_307_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_308,  flogtanh0x00000_308_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_309,  flogtanh0x00000_309_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_310,  flogtanh0x00000_310_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_311,  flogtanh0x00000_311_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_312,  flogtanh0x00000_312_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_313,  flogtanh0x00000_313_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_314,  flogtanh0x00000_314_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_315,  flogtanh0x00000_315_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_316,  flogtanh0x00000_316_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_317,  flogtanh0x00000_317_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_318,  flogtanh0x00000_318_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_319,  flogtanh0x00000_319_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_320,  flogtanh0x00000_320_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_321,  flogtanh0x00000_321_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_322,  flogtanh0x00000_322_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_323,  flogtanh0x00000_323_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_324,  flogtanh0x00000_324_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_325,  flogtanh0x00000_325_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_326,  flogtanh0x00000_326_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_327,  flogtanh0x00000_327_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_328,  flogtanh0x00000_328_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_329,  flogtanh0x00000_329_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_330,  flogtanh0x00000_330_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_331,  flogtanh0x00000_331_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_332,  flogtanh0x00000_332_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_333,  flogtanh0x00000_333_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_334,  flogtanh0x00000_334_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_335,  flogtanh0x00000_335_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_336,  flogtanh0x00000_336_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_337,  flogtanh0x00000_337_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_338,  flogtanh0x00000_338_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_339,  flogtanh0x00000_339_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_340,  flogtanh0x00000_340_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_341,  flogtanh0x00000_341_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_342,  flogtanh0x00000_342_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_343,  flogtanh0x00000_343_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_344,  flogtanh0x00000_344_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_345,  flogtanh0x00000_345_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_346,  flogtanh0x00000_346_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_347,  flogtanh0x00000_347_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_348,  flogtanh0x00000_348_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_349,  flogtanh0x00000_349_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_350,  flogtanh0x00000_350_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_351,  flogtanh0x00000_351_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_352,  flogtanh0x00000_352_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_353,  flogtanh0x00000_353_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_354,  flogtanh0x00000_354_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00000_355,  flogtanh0x00000_355_q;
wire start_d_flogtanh0x00000;
reg start_d_flogtanh0x00000_q;
always_comb begin
 flogtanh0x00000_0_q = flogtanh0x00000_0;
 flogtanh0x00000_1_q = flogtanh0x00000_1;
 flogtanh0x00000_2_q = flogtanh0x00000_2;
 flogtanh0x00000_3_q = flogtanh0x00000_3;
 flogtanh0x00000_4_q = flogtanh0x00000_4;
 flogtanh0x00000_5_q = flogtanh0x00000_5;
 flogtanh0x00000_6_q = flogtanh0x00000_6;
 flogtanh0x00000_7_q = flogtanh0x00000_7;
 flogtanh0x00000_8_q = flogtanh0x00000_8;
 flogtanh0x00000_9_q = flogtanh0x00000_9;
 flogtanh0x00000_10_q = flogtanh0x00000_10;
 flogtanh0x00000_11_q = flogtanh0x00000_11;
 flogtanh0x00000_12_q = flogtanh0x00000_12;
 flogtanh0x00000_13_q = flogtanh0x00000_13;
 flogtanh0x00000_14_q = flogtanh0x00000_14;
 flogtanh0x00000_15_q = flogtanh0x00000_15;
 flogtanh0x00000_16_q = flogtanh0x00000_16;
 flogtanh0x00000_17_q = flogtanh0x00000_17;
 flogtanh0x00000_18_q = flogtanh0x00000_18;
 flogtanh0x00000_19_q = flogtanh0x00000_19;
 flogtanh0x00000_20_q = flogtanh0x00000_20;
 flogtanh0x00000_21_q = flogtanh0x00000_21;
 flogtanh0x00000_22_q = flogtanh0x00000_22;
 flogtanh0x00000_23_q = flogtanh0x00000_23;
 flogtanh0x00000_24_q = flogtanh0x00000_24;
 flogtanh0x00000_25_q = flogtanh0x00000_25;
 flogtanh0x00000_26_q = flogtanh0x00000_26;
 flogtanh0x00000_27_q = flogtanh0x00000_27;
 flogtanh0x00000_28_q = flogtanh0x00000_28;
 flogtanh0x00000_29_q = flogtanh0x00000_29;
 flogtanh0x00000_30_q = flogtanh0x00000_30;
 flogtanh0x00000_31_q = flogtanh0x00000_31;
 flogtanh0x00000_32_q = flogtanh0x00000_32;
 flogtanh0x00000_33_q = flogtanh0x00000_33;
 flogtanh0x00000_34_q = flogtanh0x00000_34;
 flogtanh0x00000_35_q = flogtanh0x00000_35;
 flogtanh0x00000_36_q = flogtanh0x00000_36;
 flogtanh0x00000_37_q = flogtanh0x00000_37;
 flogtanh0x00000_38_q = flogtanh0x00000_38;
 flogtanh0x00000_39_q = flogtanh0x00000_39;
 flogtanh0x00000_40_q = flogtanh0x00000_40;
 flogtanh0x00000_41_q = flogtanh0x00000_41;
 flogtanh0x00000_42_q = flogtanh0x00000_42;
 flogtanh0x00000_43_q = flogtanh0x00000_43;
 flogtanh0x00000_44_q = flogtanh0x00000_44;
 flogtanh0x00000_45_q = flogtanh0x00000_45;
 flogtanh0x00000_46_q = flogtanh0x00000_46;
 flogtanh0x00000_47_q = flogtanh0x00000_47;
 flogtanh0x00000_48_q = flogtanh0x00000_48;
 flogtanh0x00000_49_q = flogtanh0x00000_49;
 flogtanh0x00000_50_q = flogtanh0x00000_50;
 flogtanh0x00000_51_q = flogtanh0x00000_51;
 flogtanh0x00000_52_q = flogtanh0x00000_52;
 flogtanh0x00000_53_q = flogtanh0x00000_53;
 flogtanh0x00000_54_q = flogtanh0x00000_54;
 flogtanh0x00000_55_q = flogtanh0x00000_55;
 flogtanh0x00000_56_q = flogtanh0x00000_56;
 flogtanh0x00000_57_q = flogtanh0x00000_57;
 flogtanh0x00000_58_q = flogtanh0x00000_58;
 flogtanh0x00000_59_q = flogtanh0x00000_59;
 flogtanh0x00000_60_q = flogtanh0x00000_60;
 flogtanh0x00000_61_q = flogtanh0x00000_61;
 flogtanh0x00000_62_q = flogtanh0x00000_62;
 flogtanh0x00000_63_q = flogtanh0x00000_63;
 flogtanh0x00000_64_q = flogtanh0x00000_64;
 flogtanh0x00000_65_q = flogtanh0x00000_65;
 flogtanh0x00000_66_q = flogtanh0x00000_66;
 flogtanh0x00000_67_q = flogtanh0x00000_67;
 flogtanh0x00000_68_q = flogtanh0x00000_68;
 flogtanh0x00000_69_q = flogtanh0x00000_69;
 flogtanh0x00000_70_q = flogtanh0x00000_70;
 flogtanh0x00000_71_q = flogtanh0x00000_71;
 flogtanh0x00000_72_q = flogtanh0x00000_72;
 flogtanh0x00000_73_q = flogtanh0x00000_73;
 flogtanh0x00000_74_q = flogtanh0x00000_74;
 flogtanh0x00000_75_q = flogtanh0x00000_75;
 flogtanh0x00000_76_q = flogtanh0x00000_76;
 flogtanh0x00000_77_q = flogtanh0x00000_77;
 flogtanh0x00000_78_q = flogtanh0x00000_78;
 flogtanh0x00000_79_q = flogtanh0x00000_79;
 flogtanh0x00000_80_q = flogtanh0x00000_80;
 flogtanh0x00000_81_q = flogtanh0x00000_81;
 flogtanh0x00000_82_q = flogtanh0x00000_82;
 flogtanh0x00000_83_q = flogtanh0x00000_83;
 flogtanh0x00000_84_q = flogtanh0x00000_84;
 flogtanh0x00000_85_q = flogtanh0x00000_85;
 flogtanh0x00000_86_q = flogtanh0x00000_86;
 flogtanh0x00000_87_q = flogtanh0x00000_87;
 flogtanh0x00000_88_q = flogtanh0x00000_88;
 flogtanh0x00000_89_q = flogtanh0x00000_89;
 flogtanh0x00000_90_q = flogtanh0x00000_90;
 flogtanh0x00000_91_q = flogtanh0x00000_91;
 flogtanh0x00000_92_q = flogtanh0x00000_92;
 flogtanh0x00000_93_q = flogtanh0x00000_93;
 flogtanh0x00000_94_q = flogtanh0x00000_94;
 flogtanh0x00000_95_q = flogtanh0x00000_95;
 flogtanh0x00000_96_q = flogtanh0x00000_96;
 flogtanh0x00000_97_q = flogtanh0x00000_97;
 flogtanh0x00000_98_q = flogtanh0x00000_98;
 flogtanh0x00000_99_q = flogtanh0x00000_99;
 flogtanh0x00000_100_q = flogtanh0x00000_100;
 flogtanh0x00000_101_q = flogtanh0x00000_101;
 flogtanh0x00000_102_q = flogtanh0x00000_102;
 flogtanh0x00000_103_q = flogtanh0x00000_103;
 flogtanh0x00000_104_q = flogtanh0x00000_104;
 flogtanh0x00000_105_q = flogtanh0x00000_105;
 flogtanh0x00000_106_q = flogtanh0x00000_106;
 flogtanh0x00000_107_q = flogtanh0x00000_107;
 flogtanh0x00000_108_q = flogtanh0x00000_108;
 flogtanh0x00000_109_q = flogtanh0x00000_109;
 flogtanh0x00000_110_q = flogtanh0x00000_110;
 flogtanh0x00000_111_q = flogtanh0x00000_111;
 flogtanh0x00000_112_q = flogtanh0x00000_112;
 flogtanh0x00000_113_q = flogtanh0x00000_113;
 flogtanh0x00000_114_q = flogtanh0x00000_114;
 flogtanh0x00000_115_q = flogtanh0x00000_115;
 flogtanh0x00000_116_q = flogtanh0x00000_116;
 flogtanh0x00000_117_q = flogtanh0x00000_117;
 flogtanh0x00000_118_q = flogtanh0x00000_118;
 flogtanh0x00000_119_q = flogtanh0x00000_119;
 flogtanh0x00000_120_q = flogtanh0x00000_120;
 flogtanh0x00000_121_q = flogtanh0x00000_121;
 flogtanh0x00000_122_q = flogtanh0x00000_122;
 flogtanh0x00000_123_q = flogtanh0x00000_123;
 flogtanh0x00000_124_q = flogtanh0x00000_124;
 flogtanh0x00000_125_q = flogtanh0x00000_125;
 flogtanh0x00000_126_q = flogtanh0x00000_126;
 flogtanh0x00000_127_q = flogtanh0x00000_127;
 flogtanh0x00000_128_q = flogtanh0x00000_128;
 flogtanh0x00000_129_q = flogtanh0x00000_129;
 flogtanh0x00000_130_q = flogtanh0x00000_130;
 flogtanh0x00000_131_q = flogtanh0x00000_131;
 flogtanh0x00000_132_q = flogtanh0x00000_132;
 flogtanh0x00000_133_q = flogtanh0x00000_133;
 flogtanh0x00000_134_q = flogtanh0x00000_134;
 flogtanh0x00000_135_q = flogtanh0x00000_135;
 flogtanh0x00000_136_q = flogtanh0x00000_136;
 flogtanh0x00000_137_q = flogtanh0x00000_137;
 flogtanh0x00000_138_q = flogtanh0x00000_138;
 flogtanh0x00000_139_q = flogtanh0x00000_139;
 flogtanh0x00000_140_q = flogtanh0x00000_140;
 flogtanh0x00000_141_q = flogtanh0x00000_141;
 flogtanh0x00000_142_q = flogtanh0x00000_142;
 flogtanh0x00000_143_q = flogtanh0x00000_143;
 flogtanh0x00000_144_q = flogtanh0x00000_144;
 flogtanh0x00000_145_q = flogtanh0x00000_145;
 flogtanh0x00000_146_q = flogtanh0x00000_146;
 flogtanh0x00000_147_q = flogtanh0x00000_147;
 flogtanh0x00000_148_q = flogtanh0x00000_148;
 flogtanh0x00000_149_q = flogtanh0x00000_149;
 flogtanh0x00000_150_q = flogtanh0x00000_150;
 flogtanh0x00000_151_q = flogtanh0x00000_151;
 flogtanh0x00000_152_q = flogtanh0x00000_152;
 flogtanh0x00000_153_q = flogtanh0x00000_153;
 flogtanh0x00000_154_q = flogtanh0x00000_154;
 flogtanh0x00000_155_q = flogtanh0x00000_155;
 flogtanh0x00000_156_q = flogtanh0x00000_156;
 flogtanh0x00000_157_q = flogtanh0x00000_157;
 flogtanh0x00000_158_q = flogtanh0x00000_158;
 flogtanh0x00000_159_q = flogtanh0x00000_159;
 flogtanh0x00000_160_q = flogtanh0x00000_160;
 flogtanh0x00000_161_q = flogtanh0x00000_161;
 flogtanh0x00000_162_q = flogtanh0x00000_162;
 flogtanh0x00000_163_q = flogtanh0x00000_163;
 flogtanh0x00000_164_q = flogtanh0x00000_164;
 flogtanh0x00000_165_q = flogtanh0x00000_165;
 flogtanh0x00000_166_q = flogtanh0x00000_166;
 flogtanh0x00000_167_q = flogtanh0x00000_167;
 flogtanh0x00000_168_q = flogtanh0x00000_168;
 flogtanh0x00000_169_q = flogtanh0x00000_169;
 flogtanh0x00000_170_q = flogtanh0x00000_170;
 flogtanh0x00000_171_q = flogtanh0x00000_171;
 flogtanh0x00000_172_q = flogtanh0x00000_172;
 flogtanh0x00000_173_q = flogtanh0x00000_173;
 flogtanh0x00000_174_q = flogtanh0x00000_174;
 flogtanh0x00000_175_q = flogtanh0x00000_175;
 flogtanh0x00000_176_q = flogtanh0x00000_176;
 flogtanh0x00000_177_q = flogtanh0x00000_177;
 flogtanh0x00000_178_q = flogtanh0x00000_178;
 flogtanh0x00000_179_q = flogtanh0x00000_179;
 flogtanh0x00000_180_q = flogtanh0x00000_180;
 flogtanh0x00000_181_q = flogtanh0x00000_181;
 flogtanh0x00000_182_q = flogtanh0x00000_182;
 flogtanh0x00000_183_q = flogtanh0x00000_183;
 flogtanh0x00000_184_q = flogtanh0x00000_184;
 flogtanh0x00000_185_q = flogtanh0x00000_185;
 flogtanh0x00000_186_q = flogtanh0x00000_186;
 flogtanh0x00000_187_q = flogtanh0x00000_187;
 flogtanh0x00000_188_q = flogtanh0x00000_188;
 flogtanh0x00000_189_q = flogtanh0x00000_189;
 flogtanh0x00000_190_q = flogtanh0x00000_190;
 flogtanh0x00000_191_q = flogtanh0x00000_191;
 flogtanh0x00000_192_q = flogtanh0x00000_192;
 flogtanh0x00000_193_q = flogtanh0x00000_193;
 flogtanh0x00000_194_q = flogtanh0x00000_194;
 flogtanh0x00000_195_q = flogtanh0x00000_195;
 flogtanh0x00000_196_q = flogtanh0x00000_196;
 flogtanh0x00000_197_q = flogtanh0x00000_197;
 flogtanh0x00000_198_q = flogtanh0x00000_198;
 flogtanh0x00000_199_q = flogtanh0x00000_199;
 flogtanh0x00000_200_q = flogtanh0x00000_200;
 flogtanh0x00000_201_q = flogtanh0x00000_201;
 flogtanh0x00000_202_q = flogtanh0x00000_202;
 flogtanh0x00000_203_q = flogtanh0x00000_203;
 flogtanh0x00000_204_q = flogtanh0x00000_204;
 flogtanh0x00000_205_q = flogtanh0x00000_205;
 flogtanh0x00000_206_q = flogtanh0x00000_206;
 flogtanh0x00000_207_q = flogtanh0x00000_207;
 flogtanh0x00000_208_q = flogtanh0x00000_208;
 flogtanh0x00000_209_q = flogtanh0x00000_209;
 flogtanh0x00000_210_q = flogtanh0x00000_210;
 flogtanh0x00000_211_q = flogtanh0x00000_211;
 flogtanh0x00000_212_q = flogtanh0x00000_212;
 flogtanh0x00000_213_q = flogtanh0x00000_213;
 flogtanh0x00000_214_q = flogtanh0x00000_214;
 flogtanh0x00000_215_q = flogtanh0x00000_215;
 flogtanh0x00000_216_q = flogtanh0x00000_216;
 flogtanh0x00000_217_q = flogtanh0x00000_217;
 flogtanh0x00000_218_q = flogtanh0x00000_218;
 flogtanh0x00000_219_q = flogtanh0x00000_219;
 flogtanh0x00000_220_q = flogtanh0x00000_220;
 flogtanh0x00000_221_q = flogtanh0x00000_221;
 flogtanh0x00000_222_q = flogtanh0x00000_222;
 flogtanh0x00000_223_q = flogtanh0x00000_223;
 flogtanh0x00000_224_q = flogtanh0x00000_224;
 flogtanh0x00000_225_q = flogtanh0x00000_225;
 flogtanh0x00000_226_q = flogtanh0x00000_226;
 flogtanh0x00000_227_q = flogtanh0x00000_227;
 flogtanh0x00000_228_q = flogtanh0x00000_228;
 flogtanh0x00000_229_q = flogtanh0x00000_229;
 flogtanh0x00000_230_q = flogtanh0x00000_230;
 flogtanh0x00000_231_q = flogtanh0x00000_231;
 flogtanh0x00000_232_q = flogtanh0x00000_232;
 flogtanh0x00000_233_q = flogtanh0x00000_233;
 flogtanh0x00000_234_q = flogtanh0x00000_234;
 flogtanh0x00000_235_q = flogtanh0x00000_235;
 flogtanh0x00000_236_q = flogtanh0x00000_236;
 flogtanh0x00000_237_q = flogtanh0x00000_237;
 flogtanh0x00000_238_q = flogtanh0x00000_238;
 flogtanh0x00000_239_q = flogtanh0x00000_239;
 flogtanh0x00000_240_q = flogtanh0x00000_240;
 flogtanh0x00000_241_q = flogtanh0x00000_241;
 flogtanh0x00000_242_q = flogtanh0x00000_242;
 flogtanh0x00000_243_q = flogtanh0x00000_243;
 flogtanh0x00000_244_q = flogtanh0x00000_244;
 flogtanh0x00000_245_q = flogtanh0x00000_245;
 flogtanh0x00000_246_q = flogtanh0x00000_246;
 flogtanh0x00000_247_q = flogtanh0x00000_247;
 flogtanh0x00000_248_q = flogtanh0x00000_248;
 flogtanh0x00000_249_q = flogtanh0x00000_249;
 flogtanh0x00000_250_q = flogtanh0x00000_250;
 flogtanh0x00000_251_q = flogtanh0x00000_251;
 flogtanh0x00000_252_q = flogtanh0x00000_252;
 flogtanh0x00000_253_q = flogtanh0x00000_253;
 flogtanh0x00000_254_q = flogtanh0x00000_254;
 flogtanh0x00000_255_q = flogtanh0x00000_255;
 flogtanh0x00000_256_q = flogtanh0x00000_256;
 flogtanh0x00000_257_q = flogtanh0x00000_257;
 flogtanh0x00000_258_q = flogtanh0x00000_258;
 flogtanh0x00000_259_q = flogtanh0x00000_259;
 flogtanh0x00000_260_q = flogtanh0x00000_260;
 flogtanh0x00000_261_q = flogtanh0x00000_261;
 flogtanh0x00000_262_q = flogtanh0x00000_262;
 flogtanh0x00000_263_q = flogtanh0x00000_263;
 flogtanh0x00000_264_q = flogtanh0x00000_264;
 flogtanh0x00000_265_q = flogtanh0x00000_265;
 flogtanh0x00000_266_q = flogtanh0x00000_266;
 flogtanh0x00000_267_q = flogtanh0x00000_267;
 flogtanh0x00000_268_q = flogtanh0x00000_268;
 flogtanh0x00000_269_q = flogtanh0x00000_269;
 flogtanh0x00000_270_q = flogtanh0x00000_270;
 flogtanh0x00000_271_q = flogtanh0x00000_271;
 flogtanh0x00000_272_q = flogtanh0x00000_272;
 flogtanh0x00000_273_q = flogtanh0x00000_273;
 flogtanh0x00000_274_q = flogtanh0x00000_274;
 flogtanh0x00000_275_q = flogtanh0x00000_275;
 flogtanh0x00000_276_q = flogtanh0x00000_276;
 flogtanh0x00000_277_q = flogtanh0x00000_277;
 flogtanh0x00000_278_q = flogtanh0x00000_278;
 flogtanh0x00000_279_q = flogtanh0x00000_279;
 flogtanh0x00000_280_q = flogtanh0x00000_280;
 flogtanh0x00000_281_q = flogtanh0x00000_281;
 flogtanh0x00000_282_q = flogtanh0x00000_282;
 flogtanh0x00000_283_q = flogtanh0x00000_283;
 flogtanh0x00000_284_q = flogtanh0x00000_284;
 flogtanh0x00000_285_q = flogtanh0x00000_285;
 flogtanh0x00000_286_q = flogtanh0x00000_286;
 flogtanh0x00000_287_q = flogtanh0x00000_287;
 flogtanh0x00000_288_q = flogtanh0x00000_288;
 flogtanh0x00000_289_q = flogtanh0x00000_289;
 flogtanh0x00000_290_q = flogtanh0x00000_290;
 flogtanh0x00000_291_q = flogtanh0x00000_291;
 flogtanh0x00000_292_q = flogtanh0x00000_292;
 flogtanh0x00000_293_q = flogtanh0x00000_293;
 flogtanh0x00000_294_q = flogtanh0x00000_294;
 flogtanh0x00000_295_q = flogtanh0x00000_295;
 flogtanh0x00000_296_q = flogtanh0x00000_296;
 flogtanh0x00000_297_q = flogtanh0x00000_297;
 flogtanh0x00000_298_q = flogtanh0x00000_298;
 flogtanh0x00000_299_q = flogtanh0x00000_299;
 flogtanh0x00000_300_q = flogtanh0x00000_300;
 flogtanh0x00000_301_q = flogtanh0x00000_301;
 flogtanh0x00000_302_q = flogtanh0x00000_302;
 flogtanh0x00000_303_q = flogtanh0x00000_303;
 flogtanh0x00000_304_q = flogtanh0x00000_304;
 flogtanh0x00000_305_q = flogtanh0x00000_305;
 flogtanh0x00000_306_q = flogtanh0x00000_306;
 flogtanh0x00000_307_q = flogtanh0x00000_307;
 flogtanh0x00000_308_q = flogtanh0x00000_308;
 flogtanh0x00000_309_q = flogtanh0x00000_309;
 flogtanh0x00000_310_q = flogtanh0x00000_310;
 flogtanh0x00000_311_q = flogtanh0x00000_311;
 flogtanh0x00000_312_q = flogtanh0x00000_312;
 flogtanh0x00000_313_q = flogtanh0x00000_313;
 flogtanh0x00000_314_q = flogtanh0x00000_314;
 flogtanh0x00000_315_q = flogtanh0x00000_315;
 flogtanh0x00000_316_q = flogtanh0x00000_316;
 flogtanh0x00000_317_q = flogtanh0x00000_317;
 flogtanh0x00000_318_q = flogtanh0x00000_318;
 flogtanh0x00000_319_q = flogtanh0x00000_319;
 flogtanh0x00000_320_q = flogtanh0x00000_320;
 flogtanh0x00000_321_q = flogtanh0x00000_321;
 flogtanh0x00000_322_q = flogtanh0x00000_322;
 flogtanh0x00000_323_q = flogtanh0x00000_323;
 flogtanh0x00000_324_q = flogtanh0x00000_324;
 flogtanh0x00000_325_q = flogtanh0x00000_325;
 flogtanh0x00000_326_q = flogtanh0x00000_326;
 flogtanh0x00000_327_q = flogtanh0x00000_327;
 flogtanh0x00000_328_q = flogtanh0x00000_328;
 flogtanh0x00000_329_q = flogtanh0x00000_329;
 flogtanh0x00000_330_q = flogtanh0x00000_330;
 flogtanh0x00000_331_q = flogtanh0x00000_331;
 flogtanh0x00000_332_q = flogtanh0x00000_332;
 flogtanh0x00000_333_q = flogtanh0x00000_333;
 flogtanh0x00000_334_q = flogtanh0x00000_334;
 flogtanh0x00000_335_q = flogtanh0x00000_335;
 flogtanh0x00000_336_q = flogtanh0x00000_336;
 flogtanh0x00000_337_q = flogtanh0x00000_337;
 flogtanh0x00000_338_q = flogtanh0x00000_338;
 flogtanh0x00000_339_q = flogtanh0x00000_339;
 flogtanh0x00000_340_q = flogtanh0x00000_340;
 flogtanh0x00000_341_q = flogtanh0x00000_341;
 flogtanh0x00000_342_q = flogtanh0x00000_342;
 flogtanh0x00000_343_q = flogtanh0x00000_343;
 flogtanh0x00000_344_q = flogtanh0x00000_344;
 flogtanh0x00000_345_q = flogtanh0x00000_345;
 flogtanh0x00000_346_q = flogtanh0x00000_346;
 flogtanh0x00000_347_q = flogtanh0x00000_347;
 flogtanh0x00000_348_q = flogtanh0x00000_348;
 flogtanh0x00000_349_q = flogtanh0x00000_349;
 flogtanh0x00000_350_q = flogtanh0x00000_350;
 flogtanh0x00000_351_q = flogtanh0x00000_351;
 flogtanh0x00000_352_q = flogtanh0x00000_352;
 flogtanh0x00000_353_q = flogtanh0x00000_353;
 flogtanh0x00000_354_q = flogtanh0x00000_354;
 flogtanh0x00000_355_q = flogtanh0x00000_355;
 start_d_flogtanh0x00000_q =  start_d_flogtanh0x00000;
end
