reg [fgallag_WDTH -1:0] fgallag0x00006_0, fgallag0x00006_0_q;
reg [fgallag_WDTH -1:0] fgallag0x00006_1, fgallag0x00006_1_q;
reg [fgallag_WDTH -1:0] fgallag0x00006_2, fgallag0x00006_2_q;
reg [fgallag_WDTH -1:0] fgallag0x00006_3, fgallag0x00006_3_q;
reg [fgallag_WDTH -1:0] fgallag0x00006_4, fgallag0x00006_4_q;
reg [fgallag_WDTH -1:0] fgallag0x00006_5, fgallag0x00006_5_q;
reg start_d_fgallag0x00006_q ;
always_comb begin
 fgallag0x00006_0_q =  fgallag0x00006_0;
 fgallag0x00006_1_q =  fgallag0x00006_1;
 fgallag0x00006_2_q =  fgallag0x00006_2;
 fgallag0x00006_3_q =  fgallag0x00006_3;
 fgallag0x00006_4_q =  fgallag0x00006_4;
 fgallag0x00006_5_q =  fgallag0x00006_5;
 start_d_fgallag0x00006_q =  start_d_fgallag0x00005_q;
end
