              fgallag0x00002_0 = 
          (!fgallag_sel[1]) ? 
                       fgallag0x00001_0_q: 
                       fgallag0x00001_1_q;
              fgallag0x00002_1 = 
          (!fgallag_sel[1]) ? 
                       fgallag0x00001_2_q: 
                       fgallag0x00001_3_q;
              fgallag0x00002_2 = 
          (!fgallag_sel[1]) ? 
                       fgallag0x00001_4_q: 
                       fgallag0x00001_5_q;
              fgallag0x00002_3 = 
          (!fgallag_sel[1]) ? 
                       fgallag0x00001_6_q: 
                       fgallag0x00001_7_q;
              fgallag0x00002_4 = 
          (!fgallag_sel[1]) ? 
                       fgallag0x00001_8_q: 
                       fgallag0x00001_9_q;
              fgallag0x00002_5 = 
          (!fgallag_sel[1]) ? 
                       fgallag0x00001_10_q: 
                       fgallag0x00001_11_q;
              fgallag0x00002_6 = 
          (!fgallag_sel[1]) ? 
                       fgallag0x00001_12_q: 
                       fgallag0x00001_13_q;
              fgallag0x00002_7 = 
          (!fgallag_sel[1]) ? 
                       fgallag0x00001_14_q: 
                       fgallag0x00001_15_q;
              fgallag0x00002_8 = 
          (!fgallag_sel[1]) ? 
                       fgallag0x00001_16_q: 
                       fgallag0x00001_17_q;
              fgallag0x00002_9 = 
          (!fgallag_sel[1]) ? 
                       fgallag0x00001_18_q: 
                       fgallag0x00001_19_q;
              fgallag0x00002_10 = 
          (!fgallag_sel[1]) ? 
                       fgallag0x00001_20_q: 
                       fgallag0x00001_21_q;
              fgallag0x00002_11 = 
          (!fgallag_sel[1]) ? 
                       fgallag0x00001_22_q: 
                       fgallag0x00001_23_q;
              fgallag0x00002_12 = 
          (!fgallag_sel[1]) ? 
                       fgallag0x00001_24_q: 
                       fgallag0x00001_25_q;
              fgallag0x00002_13 = 
          (!fgallag_sel[1]) ? 
                       fgallag0x00001_26_q: 
                       fgallag0x00001_27_q;
              fgallag0x00002_14 = 
          (!fgallag_sel[1]) ? 
                       fgallag0x00001_28_q: 
                       fgallag0x00001_29_q;
              fgallag0x00002_15 = 
          (!fgallag_sel[1]) ? 
                       fgallag0x00001_30_q: 
                       fgallag0x00001_31_q;
              fgallag0x00002_16 = 
          (!fgallag_sel[1]) ? 
                       fgallag0x00001_32_q: 
                       fgallag0x00001_33_q;
              fgallag0x00002_17 = 
          (!fgallag_sel[1]) ? 
                       fgallag0x00001_34_q: 
                       fgallag0x00001_35_q;
              fgallag0x00002_18 = 
          (!fgallag_sel[1]) ? 
                       fgallag0x00001_36_q: 
                       fgallag0x00001_37_q;
              fgallag0x00002_19 = 
          (!fgallag_sel[1]) ? 
                       fgallag0x00001_38_q: 
                       fgallag0x00001_39_q;
              fgallag0x00002_20 = 
          (!fgallag_sel[1]) ? 
                       fgallag0x00001_40_q: 
                       fgallag0x00001_41_q;
              fgallag0x00002_21 = 
          (!fgallag_sel[1]) ? 
                       fgallag0x00001_42_q: 
                       fgallag0x00001_43_q;
              fgallag0x00002_22 = 
          (!fgallag_sel[1]) ? 
                       fgallag0x00001_44_q: 
                       fgallag0x00001_45_q;
              fgallag0x00002_23 = 
          (!fgallag_sel[1]) ? 
                       fgallag0x00001_46_q: 
                       fgallag0x00001_47_q;
              fgallag0x00002_24 = 
          (!fgallag_sel[1]) ? 
                       fgallag0x00001_48_q: 
                       fgallag0x00001_49_q;
              fgallag0x00002_25 = 
          (!fgallag_sel[1]) ? 
                       fgallag0x00001_50_q: 
                       fgallag0x00001_51_q;
              fgallag0x00002_26 = 
          (!fgallag_sel[1]) ? 
                       fgallag0x00001_52_q: 
                       fgallag0x00001_53_q;
              fgallag0x00002_27 = 
          (!fgallag_sel[1]) ? 
                       fgallag0x00001_54_q: 
                       fgallag0x00001_55_q;
              fgallag0x00002_28 = 
          (!fgallag_sel[1]) ? 
                       fgallag0x00001_56_q: 
                       fgallag0x00001_57_q;
              fgallag0x00002_29 = 
          (!fgallag_sel[1]) ? 
                       fgallag0x00001_58_q: 
                       fgallag0x00001_59_q;
              fgallag0x00002_30 = 
          (!fgallag_sel[1]) ? 
                       fgallag0x00001_60_q: 
                       fgallag0x00001_61_q;
              fgallag0x00002_31 = 
          (!fgallag_sel[1]) ? 
                       fgallag0x00001_62_q: 
                       fgallag0x00001_63_q;
              fgallag0x00002_32 = 
          (!fgallag_sel[1]) ? 
                       fgallag0x00001_64_q: 
                       fgallag0x00001_65_q;
               fgallag0x00002_33 =  fgallag0x00001_66_q ;
               fgallag0x00002_34 =  fgallag0x00001_68_q ;
               fgallag0x00002_35 =  fgallag0x00001_70_q ;
              fgallag0x00002_36 = 
          (!fgallag_sel[1]) ? 
                       fgallag0x00001_72_q: 
                       fgallag0x00001_73_q;
              fgallag0x00002_37 = 
          (!fgallag_sel[1]) ? 
                       fgallag0x00001_74_q: 
                       fgallag0x00001_75_q;
              fgallag0x00002_38 = 
          (!fgallag_sel[1]) ? 
                       fgallag0x00001_76_q: 
                       fgallag0x00001_77_q;
               fgallag0x00002_39 =  fgallag0x00001_78_q ;
              fgallag0x00002_40 = 
          (!fgallag_sel[1]) ? 
                       fgallag0x00001_80_q: 
                       fgallag0x00001_81_q;
              fgallag0x00002_41 = 
          (!fgallag_sel[1]) ? 
                       fgallag0x00001_82_q: 
                       fgallag0x00001_83_q;
               fgallag0x00002_42 =  fgallag0x00001_84_q ;
              fgallag0x00002_43 = 
          (!fgallag_sel[1]) ? 
                       fgallag0x00001_86_q: 
                       fgallag0x00001_87_q;
               fgallag0x00002_44 =  fgallag0x00001_88_q ;
              fgallag0x00002_45 = 
          (!fgallag_sel[1]) ? 
                       fgallag0x00001_90_q: 
                       fgallag0x00001_91_q;
               fgallag0x00002_46 =  fgallag0x00001_92_q ;
               fgallag0x00002_47 =  fgallag0x00001_94_q ;
               fgallag0x00002_48 =  fgallag0x00001_96_q ;
               fgallag0x00002_49 =  fgallag0x00001_98_q ;
              fgallag0x00002_50 = 
          (!fgallag_sel[1]) ? 
                       fgallag0x00001_100_q: 
                       fgallag0x00001_101_q;
               fgallag0x00002_51 =  fgallag0x00001_102_q ;
               fgallag0x00002_52 =  fgallag0x00001_104_q ;
              fgallag0x00002_53 = 
          (!fgallag_sel[1]) ? 
                       fgallag0x00001_106_q: 
                       fgallag0x00001_107_q;
               fgallag0x00002_54 =  fgallag0x00001_108_q ;
               fgallag0x00002_55 =  fgallag0x00001_110_q ;
               fgallag0x00002_56 =  fgallag0x00001_112_q ;
              fgallag0x00002_57 = 
          (!fgallag_sel[1]) ? 
                       fgallag0x00001_114_q: 
                       fgallag0x00001_115_q;
               fgallag0x00002_58 =  fgallag0x00001_116_q ;
               fgallag0x00002_59 =  fgallag0x00001_118_q ;
               fgallag0x00002_60 =  fgallag0x00001_120_q ;
               fgallag0x00002_61 =  fgallag0x00001_122_q ;
               fgallag0x00002_62 =  fgallag0x00001_124_q ;
              fgallag0x00002_63 = 
          (!fgallag_sel[1]) ? 
                       fgallag0x00001_126_q: 
                       fgallag0x00001_127_q;
               fgallag0x00002_64 =  fgallag0x00001_128_q ;
               fgallag0x00002_65 =  fgallag0x00001_130_q ;
               fgallag0x00002_66 =  fgallag0x00001_132_q ;
               fgallag0x00002_67 =  fgallag0x00001_134_q ;
               fgallag0x00002_68 =  fgallag0x00001_136_q ;
               fgallag0x00002_69 =  fgallag0x00001_138_q ;
               fgallag0x00002_70 =  fgallag0x00001_140_q ;
              fgallag0x00002_71 = 
          (!fgallag_sel[1]) ? 
                       fgallag0x00001_142_q: 
                       fgallag0x00001_143_q;
               fgallag0x00002_72 =  fgallag0x00001_144_q ;
               fgallag0x00002_73 =  fgallag0x00001_146_q ;
               fgallag0x00002_74 =  fgallag0x00001_148_q ;
               fgallag0x00002_75 =  fgallag0x00001_150_q ;
               fgallag0x00002_76 =  fgallag0x00001_152_q ;
               fgallag0x00002_77 =  fgallag0x00001_154_q ;
               fgallag0x00002_78 =  fgallag0x00001_156_q ;
               fgallag0x00002_79 =  fgallag0x00001_158_q ;
               fgallag0x00002_80 =  fgallag0x00001_160_q ;
               fgallag0x00002_81 =  fgallag0x00001_162_q ;
               fgallag0x00002_82 =  fgallag0x00001_164_q ;
               fgallag0x00002_83 =  fgallag0x00001_166_q ;
               fgallag0x00002_84 =  fgallag0x00001_168_q ;
               fgallag0x00002_85 =  fgallag0x00001_170_q ;
               fgallag0x00002_86 =  fgallag0x00001_172_q ;
               fgallag0x00002_87 =  fgallag0x00001_174_q ;
               fgallag0x00002_88 =  fgallag0x00001_176_q ;
               fgallag0x00002_89 =  0;
