`ifndef LDPC_CSR_VH
`define LDPC_CSR_VH
`define LDPC_CSR_LDPC_ENC_MSG_IN_0_MSG_IN_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_MSG_IN_0_MSG_IN_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_MSG_IN_0_MSG_IN_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_MSG_IN_0_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_0_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_0_BYTE_OFFSET 13'h0000
`define LDPC_CSR_LDPC_ENC_MSG_IN_1_MSG_IN_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_MSG_IN_1_MSG_IN_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_MSG_IN_1_MSG_IN_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_MSG_IN_1_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_1_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_1_BYTE_OFFSET 13'h0004
`define LDPC_CSR_LDPC_ENC_MSG_IN_2_MSG_IN_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_MSG_IN_2_MSG_IN_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_MSG_IN_2_MSG_IN_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_MSG_IN_2_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_2_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_2_BYTE_OFFSET 13'h0008
`define LDPC_CSR_LDPC_ENC_MSG_IN_3_MSG_IN_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_MSG_IN_3_MSG_IN_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_MSG_IN_3_MSG_IN_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_MSG_IN_3_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_3_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_3_BYTE_OFFSET 13'h000c
`define LDPC_CSR_LDPC_ENC_MSG_IN_4_MSG_IN_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_MSG_IN_4_MSG_IN_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_MSG_IN_4_MSG_IN_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_MSG_IN_4_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_4_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_4_BYTE_OFFSET 13'h0010
`define LDPC_CSR_LDPC_ENC_MSG_IN_5_MSG_IN_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_MSG_IN_5_MSG_IN_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_MSG_IN_5_MSG_IN_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_MSG_IN_5_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_5_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_5_BYTE_OFFSET 13'h0014
`define LDPC_CSR_LDPC_ENC_MSG_IN_6_MSG_IN_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_MSG_IN_6_MSG_IN_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_MSG_IN_6_MSG_IN_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_MSG_IN_6_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_6_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_6_BYTE_OFFSET 13'h0018
`define LDPC_CSR_LDPC_ENC_MSG_IN_7_MSG_IN_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_MSG_IN_7_MSG_IN_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_MSG_IN_7_MSG_IN_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_MSG_IN_7_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_7_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_7_BYTE_OFFSET 13'h001c
`define LDPC_CSR_LDPC_ENC_MSG_IN_8_MSG_IN_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_MSG_IN_8_MSG_IN_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_MSG_IN_8_MSG_IN_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_MSG_IN_8_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_8_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_8_BYTE_OFFSET 13'h0020
`define LDPC_CSR_LDPC_ENC_MSG_IN_9_MSG_IN_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_MSG_IN_9_MSG_IN_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_MSG_IN_9_MSG_IN_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_MSG_IN_9_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_9_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_9_BYTE_OFFSET 13'h0024
`define LDPC_CSR_LDPC_ENC_MSG_IN_10_MSG_IN_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_MSG_IN_10_MSG_IN_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_MSG_IN_10_MSG_IN_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_MSG_IN_10_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_10_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_10_BYTE_OFFSET 13'h0028
`define LDPC_CSR_LDPC_ENC_MSG_IN_11_MSG_IN_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_MSG_IN_11_MSG_IN_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_MSG_IN_11_MSG_IN_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_MSG_IN_11_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_11_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_11_BYTE_OFFSET 13'h002c
`define LDPC_CSR_LDPC_ENC_MSG_IN_12_MSG_IN_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_MSG_IN_12_MSG_IN_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_MSG_IN_12_MSG_IN_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_MSG_IN_12_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_12_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_12_BYTE_OFFSET 13'h0030
`define LDPC_CSR_LDPC_ENC_MSG_IN_13_MSG_IN_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_MSG_IN_13_MSG_IN_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_MSG_IN_13_MSG_IN_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_MSG_IN_13_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_13_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_13_BYTE_OFFSET 13'h0034
`define LDPC_CSR_LDPC_ENC_MSG_IN_14_MSG_IN_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_MSG_IN_14_MSG_IN_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_MSG_IN_14_MSG_IN_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_MSG_IN_14_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_14_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_14_BYTE_OFFSET 13'h0038
`define LDPC_CSR_LDPC_ENC_MSG_IN_15_MSG_IN_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_MSG_IN_15_MSG_IN_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_MSG_IN_15_MSG_IN_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_MSG_IN_15_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_15_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_15_BYTE_OFFSET 13'h003c
`define LDPC_CSR_LDPC_ENC_MSG_IN_16_MSG_IN_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_MSG_IN_16_MSG_IN_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_MSG_IN_16_MSG_IN_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_MSG_IN_16_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_16_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_16_BYTE_OFFSET 13'h0040
`define LDPC_CSR_LDPC_ENC_MSG_IN_17_MSG_IN_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_MSG_IN_17_MSG_IN_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_MSG_IN_17_MSG_IN_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_MSG_IN_17_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_17_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_17_BYTE_OFFSET 13'h0044
`define LDPC_CSR_LDPC_ENC_MSG_IN_18_MSG_IN_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_MSG_IN_18_MSG_IN_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_MSG_IN_18_MSG_IN_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_MSG_IN_18_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_18_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_18_BYTE_OFFSET 13'h0048
`define LDPC_CSR_LDPC_ENC_MSG_IN_19_MSG_IN_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_MSG_IN_19_MSG_IN_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_MSG_IN_19_MSG_IN_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_MSG_IN_19_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_19_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_19_BYTE_OFFSET 13'h004c
`define LDPC_CSR_LDPC_ENC_MSG_IN_20_MSG_IN_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_MSG_IN_20_MSG_IN_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_MSG_IN_20_MSG_IN_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_MSG_IN_20_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_20_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_20_BYTE_OFFSET 13'h0050
`define LDPC_CSR_LDPC_ENC_MSG_IN_21_MSG_IN_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_MSG_IN_21_MSG_IN_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_MSG_IN_21_MSG_IN_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_MSG_IN_21_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_21_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_21_BYTE_OFFSET 13'h0054
`define LDPC_CSR_LDPC_ENC_MSG_IN_22_MSG_IN_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_MSG_IN_22_MSG_IN_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_MSG_IN_22_MSG_IN_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_MSG_IN_22_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_22_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_22_BYTE_OFFSET 13'h0058
`define LDPC_CSR_LDPC_ENC_MSG_IN_23_MSG_IN_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_MSG_IN_23_MSG_IN_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_MSG_IN_23_MSG_IN_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_MSG_IN_23_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_23_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_23_BYTE_OFFSET 13'h005c
`define LDPC_CSR_LDPC_ENC_MSG_IN_24_MSG_IN_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_MSG_IN_24_MSG_IN_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_MSG_IN_24_MSG_IN_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_MSG_IN_24_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_24_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_24_BYTE_OFFSET 13'h0060
`define LDPC_CSR_LDPC_ENC_MSG_IN_25_MSG_IN_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_MSG_IN_25_MSG_IN_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_MSG_IN_25_MSG_IN_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_MSG_IN_25_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_25_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_25_BYTE_OFFSET 13'h0064
`define LDPC_CSR_LDPC_ENC_MSG_IN_26_MSG_IN_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_MSG_IN_26_MSG_IN_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_MSG_IN_26_MSG_IN_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_MSG_IN_26_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_26_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_26_BYTE_OFFSET 13'h0068
`define LDPC_CSR_LDPC_ENC_MSG_IN_27_MSG_IN_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_MSG_IN_27_MSG_IN_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_MSG_IN_27_MSG_IN_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_MSG_IN_27_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_27_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_27_BYTE_OFFSET 13'h006c
`define LDPC_CSR_LDPC_ENC_MSG_IN_28_MSG_IN_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_MSG_IN_28_MSG_IN_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_MSG_IN_28_MSG_IN_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_MSG_IN_28_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_28_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_28_BYTE_OFFSET 13'h0070
`define LDPC_CSR_LDPC_ENC_MSG_IN_29_MSG_IN_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_MSG_IN_29_MSG_IN_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_MSG_IN_29_MSG_IN_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_MSG_IN_29_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_29_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_29_BYTE_OFFSET 13'h0074
`define LDPC_CSR_LDPC_ENC_MSG_IN_30_MSG_IN_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_MSG_IN_30_MSG_IN_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_MSG_IN_30_MSG_IN_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_MSG_IN_30_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_30_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_30_BYTE_OFFSET 13'h0078
`define LDPC_CSR_LDPC_ENC_MSG_IN_31_MSG_IN_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_MSG_IN_31_MSG_IN_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_MSG_IN_31_MSG_IN_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_MSG_IN_31_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_31_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_31_BYTE_OFFSET 13'h007c
`define LDPC_CSR_LDPC_ENC_MSG_IN_32_MSG_IN_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_MSG_IN_32_MSG_IN_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_MSG_IN_32_MSG_IN_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_MSG_IN_32_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_32_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_32_BYTE_OFFSET 13'h0080
`define LDPC_CSR_LDPC_ENC_MSG_IN_33_MSG_IN_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_MSG_IN_33_MSG_IN_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_MSG_IN_33_MSG_IN_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_MSG_IN_33_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_33_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_33_BYTE_OFFSET 13'h0084
`define LDPC_CSR_LDPC_ENC_MSG_IN_34_MSG_IN_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_MSG_IN_34_MSG_IN_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_MSG_IN_34_MSG_IN_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_MSG_IN_34_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_34_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_34_BYTE_OFFSET 13'h0088
`define LDPC_CSR_LDPC_ENC_MSG_IN_35_MSG_IN_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_MSG_IN_35_MSG_IN_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_MSG_IN_35_MSG_IN_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_MSG_IN_35_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_35_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_35_BYTE_OFFSET 13'h008c
`define LDPC_CSR_LDPC_ENC_MSG_IN_36_MSG_IN_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_MSG_IN_36_MSG_IN_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_MSG_IN_36_MSG_IN_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_MSG_IN_36_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_36_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_36_BYTE_OFFSET 13'h0090
`define LDPC_CSR_LDPC_ENC_MSG_IN_37_MSG_IN_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_MSG_IN_37_MSG_IN_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_MSG_IN_37_MSG_IN_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_MSG_IN_37_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_37_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_37_BYTE_OFFSET 13'h0094
`define LDPC_CSR_LDPC_ENC_MSG_IN_38_MSG_IN_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_MSG_IN_38_MSG_IN_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_MSG_IN_38_MSG_IN_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_MSG_IN_38_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_38_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_38_BYTE_OFFSET 13'h0098
`define LDPC_CSR_LDPC_ENC_MSG_IN_39_MSG_IN_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_MSG_IN_39_MSG_IN_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_MSG_IN_39_MSG_IN_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_MSG_IN_39_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_39_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_MSG_IN_39_BYTE_OFFSET 13'h009c
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_0_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_0_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_0_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_0_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_0_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_0_BYTE_OFFSET 13'h00a0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_1_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_1_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_1_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_1_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_1_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_1_BYTE_OFFSET 13'h00a4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_2_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_2_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_2_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_2_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_2_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_2_BYTE_OFFSET 13'h00a8
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_3_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_3_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_3_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_3_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_3_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_3_BYTE_OFFSET 13'h00ac
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_4_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_4_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_4_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_4_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_4_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_4_BYTE_OFFSET 13'h00b0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_5_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_5_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_5_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_5_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_5_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_5_BYTE_OFFSET 13'h00b4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_6_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_6_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_6_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_6_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_6_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_6_BYTE_OFFSET 13'h00b8
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_7_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_7_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_7_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_7_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_7_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_7_BYTE_OFFSET 13'h00bc
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_8_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_8_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_8_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_8_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_8_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_8_BYTE_OFFSET 13'h00c0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_9_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_9_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_9_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_9_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_9_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_9_BYTE_OFFSET 13'h00c4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_10_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_10_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_10_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_10_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_10_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_10_BYTE_OFFSET 13'h00c8
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_11_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_11_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_11_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_11_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_11_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_11_BYTE_OFFSET 13'h00cc
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_12_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_12_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_12_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_12_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_12_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_12_BYTE_OFFSET 13'h00d0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_13_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_13_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_13_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_13_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_13_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_13_BYTE_OFFSET 13'h00d4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_14_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_14_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_14_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_14_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_14_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_14_BYTE_OFFSET 13'h00d8
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_15_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_15_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_15_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_15_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_15_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_15_BYTE_OFFSET 13'h00dc
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_16_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_16_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_16_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_16_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_16_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_16_BYTE_OFFSET 13'h00e0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_17_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_17_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_17_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_17_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_17_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_17_BYTE_OFFSET 13'h00e4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_18_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_18_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_18_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_18_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_18_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_18_BYTE_OFFSET 13'h00e8
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_19_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_19_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_19_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_19_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_19_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_19_BYTE_OFFSET 13'h00ec
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_20_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_20_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_20_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_20_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_20_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_20_BYTE_OFFSET 13'h00f0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_21_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_21_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_21_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_21_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_21_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_21_BYTE_OFFSET 13'h00f4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_22_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_22_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_22_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_22_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_22_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_22_BYTE_OFFSET 13'h00f8
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_23_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_23_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_23_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_23_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_23_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_23_BYTE_OFFSET 13'h00fc
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_24_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_24_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_24_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_24_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_24_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_24_BYTE_OFFSET 13'h0100
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_25_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_25_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_25_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_25_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_25_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_25_BYTE_OFFSET 13'h0104
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_26_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_26_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_26_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_26_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_26_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_26_BYTE_OFFSET 13'h0108
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_27_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_27_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_27_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_27_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_27_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_27_BYTE_OFFSET 13'h010c
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_28_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_28_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_28_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_28_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_28_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_28_BYTE_OFFSET 13'h0110
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_29_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_29_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_29_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_29_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_29_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_29_BYTE_OFFSET 13'h0114
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_30_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_30_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_30_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_30_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_30_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_30_BYTE_OFFSET 13'h0118
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_31_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_31_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_31_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_31_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_31_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_31_BYTE_OFFSET 13'h011c
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_32_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_32_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_32_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_32_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_32_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_32_BYTE_OFFSET 13'h0120
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_33_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_33_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_33_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_33_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_33_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_33_BYTE_OFFSET 13'h0124
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_34_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_34_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_34_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_34_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_34_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_34_BYTE_OFFSET 13'h0128
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_35_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_35_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_35_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_35_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_35_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_35_BYTE_OFFSET 13'h012c
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_36_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_36_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_36_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_36_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_36_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_36_BYTE_OFFSET 13'h0130
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_37_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_37_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_37_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_37_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_37_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_37_BYTE_OFFSET 13'h0134
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_38_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_38_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_38_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_38_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_38_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_38_BYTE_OFFSET 13'h0138
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_39_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_39_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_39_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_39_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_39_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_39_BYTE_OFFSET 13'h013c
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_40_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_40_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_40_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_40_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_40_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_40_BYTE_OFFSET 13'h0140
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_41_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_41_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_41_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_41_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_41_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_41_BYTE_OFFSET 13'h0144
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_42_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_42_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_42_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_42_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_42_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_42_BYTE_OFFSET 13'h0148
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_43_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_43_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_43_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_43_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_43_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_43_BYTE_OFFSET 13'h014c
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_44_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_44_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_44_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_44_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_44_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_44_BYTE_OFFSET 13'h0150
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_45_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_45_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_45_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_45_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_45_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_45_BYTE_OFFSET 13'h0154
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_46_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_46_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_46_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_46_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_46_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_46_BYTE_OFFSET 13'h0158
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_47_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_47_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_47_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_47_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_47_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_47_BYTE_OFFSET 13'h015c
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_48_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_48_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_48_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_48_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_48_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_48_BYTE_OFFSET 13'h0160
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_49_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_49_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_49_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_49_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_49_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_49_BYTE_OFFSET 13'h0164
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_50_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_50_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_50_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_50_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_50_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_50_BYTE_OFFSET 13'h0168
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_51_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_51_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_51_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_51_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_51_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_51_BYTE_OFFSET 13'h016c
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_52_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_52_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_52_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_52_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_52_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_52_BYTE_OFFSET 13'h0170
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_53_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_53_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_53_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_53_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_53_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_53_BYTE_OFFSET 13'h0174
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_54_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_54_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_54_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_54_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_54_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_54_BYTE_OFFSET 13'h0178
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_55_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_55_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_55_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_55_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_55_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_55_BYTE_OFFSET 13'h017c
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_56_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_56_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_56_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_56_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_56_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_56_BYTE_OFFSET 13'h0180
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_57_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_57_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_57_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_57_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_57_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_57_BYTE_OFFSET 13'h0184
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_58_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_58_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_58_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_58_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_58_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_58_BYTE_OFFSET 13'h0188
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_59_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_59_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_59_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_59_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_59_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_59_BYTE_OFFSET 13'h018c
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_60_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_60_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_60_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_60_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_60_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_60_BYTE_OFFSET 13'h0190
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_61_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_61_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_61_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_61_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_61_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_61_BYTE_OFFSET 13'h0194
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_62_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_62_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_62_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_62_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_62_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_62_BYTE_OFFSET 13'h0198
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_63_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_63_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_63_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_63_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_63_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_63_BYTE_OFFSET 13'h019c
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_64_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_64_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_64_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_64_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_64_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_64_BYTE_OFFSET 13'h01a0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_65_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_65_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_65_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_65_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_65_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_65_BYTE_OFFSET 13'h01a4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_66_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_66_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_66_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_66_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_66_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_66_BYTE_OFFSET 13'h01a8
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_67_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_67_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_67_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_67_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_67_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_67_BYTE_OFFSET 13'h01ac
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_68_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_68_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_68_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_68_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_68_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_68_BYTE_OFFSET 13'h01b0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_69_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_69_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_69_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_69_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_69_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_69_BYTE_OFFSET 13'h01b4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_70_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_70_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_70_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_70_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_70_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_70_BYTE_OFFSET 13'h01b8
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_71_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_71_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_71_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_71_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_71_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_71_BYTE_OFFSET 13'h01bc
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_72_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_72_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_72_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_72_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_72_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_72_BYTE_OFFSET 13'h01c0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_73_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_73_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_73_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_73_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_73_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_73_BYTE_OFFSET 13'h01c4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_74_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_74_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_74_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_74_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_74_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_74_BYTE_OFFSET 13'h01c8
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_75_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_75_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_75_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_75_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_75_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_75_BYTE_OFFSET 13'h01cc
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_76_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_76_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_76_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_76_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_76_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_76_BYTE_OFFSET 13'h01d0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_77_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_77_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_77_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_77_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_77_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_77_BYTE_OFFSET 13'h01d4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_78_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_78_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_78_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_78_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_78_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_78_BYTE_OFFSET 13'h01d8
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_79_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_79_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_79_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_79_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_79_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_79_BYTE_OFFSET 13'h01dc
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_80_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_80_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_80_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_80_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_80_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_80_BYTE_OFFSET 13'h01e0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_81_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_81_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_81_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_81_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_81_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_81_BYTE_OFFSET 13'h01e4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_82_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_82_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_82_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_82_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_82_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_82_BYTE_OFFSET 13'h01e8
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_83_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_83_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_83_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_83_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_83_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_83_BYTE_OFFSET 13'h01ec
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_84_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_84_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_84_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_84_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_84_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_84_BYTE_OFFSET 13'h01f0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_85_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_85_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_85_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_85_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_85_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_85_BYTE_OFFSET 13'h01f4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_86_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_86_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_86_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_86_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_86_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_86_BYTE_OFFSET 13'h01f8
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_87_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_87_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_87_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_87_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_87_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_87_BYTE_OFFSET 13'h01fc
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_88_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_88_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_88_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_88_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_88_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_88_BYTE_OFFSET 13'h0200
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_89_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_89_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_89_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_89_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_89_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_89_BYTE_OFFSET 13'h0204
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_90_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_90_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_90_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_90_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_90_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_90_BYTE_OFFSET 13'h0208
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_91_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_91_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_91_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_91_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_91_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_91_BYTE_OFFSET 13'h020c
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_92_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_92_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_92_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_92_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_92_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_92_BYTE_OFFSET 13'h0210
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_93_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_93_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_93_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_93_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_93_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_93_BYTE_OFFSET 13'h0214
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_94_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_94_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_94_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_94_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_94_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_94_BYTE_OFFSET 13'h0218
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_95_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_95_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_95_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_95_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_95_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_95_BYTE_OFFSET 13'h021c
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_96_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_96_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_96_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_96_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_96_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_96_BYTE_OFFSET 13'h0220
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_97_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_97_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_97_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_97_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_97_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_97_BYTE_OFFSET 13'h0224
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_98_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_98_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_98_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_98_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_98_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_98_BYTE_OFFSET 13'h0228
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_99_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_99_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_99_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_99_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_99_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_99_BYTE_OFFSET 13'h022c
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_100_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_100_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_100_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_100_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_100_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_100_BYTE_OFFSET 13'h0230
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_101_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_101_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_101_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_101_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_101_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_101_BYTE_OFFSET 13'h0234
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_102_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_102_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_102_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_102_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_102_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_102_BYTE_OFFSET 13'h0238
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_103_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_103_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_103_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_103_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_103_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_103_BYTE_OFFSET 13'h023c
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_104_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_104_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_104_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_104_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_104_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_104_BYTE_OFFSET 13'h0240
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_105_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_105_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_105_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_105_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_105_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_105_BYTE_OFFSET 13'h0244
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_106_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_106_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_106_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_106_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_106_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_106_BYTE_OFFSET 13'h0248
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_107_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_107_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_107_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_107_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_107_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_107_BYTE_OFFSET 13'h024c
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_108_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_108_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_108_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_108_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_108_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_108_BYTE_OFFSET 13'h0250
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_109_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_109_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_109_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_109_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_109_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_109_BYTE_OFFSET 13'h0254
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_110_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_110_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_110_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_110_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_110_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_110_BYTE_OFFSET 13'h0258
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_111_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_111_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_111_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_111_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_111_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_111_BYTE_OFFSET 13'h025c
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_112_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_112_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_112_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_112_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_112_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_112_BYTE_OFFSET 13'h0260
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_113_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_113_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_113_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_113_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_113_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_113_BYTE_OFFSET 13'h0264
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_114_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_114_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_114_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_114_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_114_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_114_BYTE_OFFSET 13'h0268
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_115_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_115_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_115_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_115_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_115_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_115_BYTE_OFFSET 13'h026c
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_116_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_116_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_116_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_116_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_116_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_116_BYTE_OFFSET 13'h0270
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_117_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_117_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_117_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_117_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_117_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_117_BYTE_OFFSET 13'h0274
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_118_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_118_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_118_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_118_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_118_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_118_BYTE_OFFSET 13'h0278
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_119_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_119_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_119_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_119_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_119_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_119_BYTE_OFFSET 13'h027c
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_120_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_120_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_120_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_120_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_120_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_120_BYTE_OFFSET 13'h0280
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_121_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_121_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_121_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_121_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_121_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_121_BYTE_OFFSET 13'h0284
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_122_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_122_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_122_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_122_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_122_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_122_BYTE_OFFSET 13'h0288
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_123_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_123_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_123_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_123_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_123_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_123_BYTE_OFFSET 13'h028c
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_124_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_124_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_124_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_124_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_124_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_124_BYTE_OFFSET 13'h0290
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_125_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_125_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_125_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_125_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_125_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_125_BYTE_OFFSET 13'h0294
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_126_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_126_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_126_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_126_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_126_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_126_BYTE_OFFSET 13'h0298
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_127_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_127_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_127_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_127_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_127_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_127_BYTE_OFFSET 13'h029c
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_128_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_128_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_128_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_128_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_128_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_128_BYTE_OFFSET 13'h02a0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_129_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_129_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_129_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_129_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_129_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_129_BYTE_OFFSET 13'h02a4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_130_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_130_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_130_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_130_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_130_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_130_BYTE_OFFSET 13'h02a8
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_131_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_131_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_131_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_131_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_131_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_131_BYTE_OFFSET 13'h02ac
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_132_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_132_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_132_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_132_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_132_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_132_BYTE_OFFSET 13'h02b0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_133_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_133_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_133_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_133_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_133_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_133_BYTE_OFFSET 13'h02b4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_134_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_134_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_134_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_134_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_134_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_134_BYTE_OFFSET 13'h02b8
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_135_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_135_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_135_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_135_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_135_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_135_BYTE_OFFSET 13'h02bc
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_136_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_136_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_136_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_136_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_136_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_136_BYTE_OFFSET 13'h02c0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_137_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_137_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_137_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_137_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_137_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_137_BYTE_OFFSET 13'h02c4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_138_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_138_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_138_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_138_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_138_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_138_BYTE_OFFSET 13'h02c8
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_139_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_139_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_139_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_139_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_139_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_139_BYTE_OFFSET 13'h02cc
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_140_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_140_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_140_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_140_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_140_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_140_BYTE_OFFSET 13'h02d0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_141_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_141_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_141_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_141_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_141_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_141_BYTE_OFFSET 13'h02d4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_142_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_142_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_142_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_142_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_142_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_142_BYTE_OFFSET 13'h02d8
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_143_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_143_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_143_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_143_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_143_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_143_BYTE_OFFSET 13'h02dc
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_144_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_144_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_144_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_144_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_144_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_144_BYTE_OFFSET 13'h02e0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_145_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_145_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_145_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_145_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_145_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_145_BYTE_OFFSET 13'h02e4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_146_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_146_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_146_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_146_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_146_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_146_BYTE_OFFSET 13'h02e8
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_147_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_147_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_147_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_147_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_147_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_147_BYTE_OFFSET 13'h02ec
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_148_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_148_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_148_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_148_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_148_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_148_BYTE_OFFSET 13'h02f0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_149_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_149_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_149_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_149_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_149_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_149_BYTE_OFFSET 13'h02f4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_150_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_150_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_150_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_150_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_150_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_150_BYTE_OFFSET 13'h02f8
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_151_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_151_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_151_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_151_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_151_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_151_BYTE_OFFSET 13'h02fc
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_152_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_152_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_152_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_152_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_152_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_152_BYTE_OFFSET 13'h0300
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_153_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_153_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_153_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_153_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_153_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_153_BYTE_OFFSET 13'h0304
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_154_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_154_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_154_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_154_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_154_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_154_BYTE_OFFSET 13'h0308
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_155_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_155_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_155_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_155_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_155_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_155_BYTE_OFFSET 13'h030c
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_156_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_156_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_156_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_156_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_156_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_156_BYTE_OFFSET 13'h0310
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_157_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_157_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_157_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_157_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_157_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_157_BYTE_OFFSET 13'h0314
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_158_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_158_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_158_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_158_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_158_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_158_BYTE_OFFSET 13'h0318
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_159_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_159_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_159_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_159_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_159_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_159_BYTE_OFFSET 13'h031c
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_160_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_160_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_160_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_160_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_160_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_160_BYTE_OFFSET 13'h0320
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_161_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_161_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_161_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_161_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_161_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_161_BYTE_OFFSET 13'h0324
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_162_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_162_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_162_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_162_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_162_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_162_BYTE_OFFSET 13'h0328
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_163_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_163_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_163_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_163_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_163_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_163_BYTE_OFFSET 13'h032c
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_164_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_164_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_164_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_164_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_164_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_164_BYTE_OFFSET 13'h0330
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_165_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_165_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_165_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_165_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_165_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_165_BYTE_OFFSET 13'h0334
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_166_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_166_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_166_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_166_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_166_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_166_BYTE_OFFSET 13'h0338
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_167_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_167_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_167_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_167_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_167_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_167_BYTE_OFFSET 13'h033c
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_168_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_168_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_168_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_168_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_168_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_168_BYTE_OFFSET 13'h0340
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_169_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_169_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_169_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_169_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_169_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_169_BYTE_OFFSET 13'h0344
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_170_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_170_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_170_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_170_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_170_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_170_BYTE_OFFSET 13'h0348
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_171_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_171_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_171_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_171_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_171_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_171_BYTE_OFFSET 13'h034c
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_172_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_172_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_172_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_172_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_172_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_172_BYTE_OFFSET 13'h0350
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_173_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_173_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_173_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_173_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_173_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_173_BYTE_OFFSET 13'h0354
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_174_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_174_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_174_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_174_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_174_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_174_BYTE_OFFSET 13'h0358
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_175_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_175_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_175_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_175_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_175_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_175_BYTE_OFFSET 13'h035c
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_176_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_176_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_176_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_176_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_176_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_176_BYTE_OFFSET 13'h0360
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_177_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_177_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_177_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_177_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_177_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_177_BYTE_OFFSET 13'h0364
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_178_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_178_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_178_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_178_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_178_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_178_BYTE_OFFSET 13'h0368
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_179_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_179_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_179_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_179_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_179_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_179_BYTE_OFFSET 13'h036c
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_180_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_180_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_180_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_180_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_180_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_180_BYTE_OFFSET 13'h0370
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_181_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_181_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_181_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_181_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_181_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_181_BYTE_OFFSET 13'h0374
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_182_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_182_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_182_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_182_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_182_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_182_BYTE_OFFSET 13'h0378
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_183_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_183_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_183_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_183_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_183_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_183_BYTE_OFFSET 13'h037c
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_184_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_184_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_184_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_184_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_184_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_184_BYTE_OFFSET 13'h0380
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_185_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_185_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_185_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_185_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_185_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_185_BYTE_OFFSET 13'h0384
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_186_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_186_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_186_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_186_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_186_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_186_BYTE_OFFSET 13'h0388
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_187_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_187_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_187_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_187_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_187_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_187_BYTE_OFFSET 13'h038c
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_188_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_188_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_188_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_188_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_188_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_188_BYTE_OFFSET 13'h0390
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_189_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_189_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_189_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_189_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_189_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_189_BYTE_OFFSET 13'h0394
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_190_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_190_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_190_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_190_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_190_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_190_BYTE_OFFSET 13'h0398
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_191_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_191_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_191_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_191_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_191_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_191_BYTE_OFFSET 13'h039c
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_192_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_192_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_192_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_192_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_192_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_192_BYTE_OFFSET 13'h03a0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_193_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_193_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_193_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_193_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_193_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_193_BYTE_OFFSET 13'h03a4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_194_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_194_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_194_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_194_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_194_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_194_BYTE_OFFSET 13'h03a8
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_195_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_195_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_195_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_195_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_195_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_195_BYTE_OFFSET 13'h03ac
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_196_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_196_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_196_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_196_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_196_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_196_BYTE_OFFSET 13'h03b0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_197_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_197_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_197_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_197_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_197_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_197_BYTE_OFFSET 13'h03b4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_198_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_198_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_198_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_198_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_198_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_198_BYTE_OFFSET 13'h03b8
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_199_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_199_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_199_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_199_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_199_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_199_BYTE_OFFSET 13'h03bc
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_200_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_200_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_200_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_200_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_200_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_200_BYTE_OFFSET 13'h03c0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_201_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_201_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_201_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_201_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_201_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_201_BYTE_OFFSET 13'h03c4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_202_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_202_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_202_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_202_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_202_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_202_BYTE_OFFSET 13'h03c8
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_203_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_203_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_203_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_203_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_203_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_203_BYTE_OFFSET 13'h03cc
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_204_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_204_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_204_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_204_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_204_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_204_BYTE_OFFSET 13'h03d0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_205_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_205_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_205_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_205_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_205_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_205_BYTE_OFFSET 13'h03d4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_206_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_206_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_206_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_206_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_206_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_206_BYTE_OFFSET 13'h03d8
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_207_ENC_CODEWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_207_ENC_CODEWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_207_ENC_CODEWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_207_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_207_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_OUT_207_BYTE_OFFSET 13'h03dc
`define LDPC_CSR_LDPC_ENC_CODEWRD_VLD_ENC_CODEWORD_VALID_BIT_WIDTH 1
`define LDPC_CSR_LDPC_ENC_CODEWRD_VLD_ENC_CODEWORD_VALID_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_ENC_CODEWRD_VLD_ENC_CODEWORD_VALID_BIT_OFFSET 0
`define LDPC_CSR_LDPC_ENC_CODEWRD_VLD_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_VLD_BYTE_SIZE 4
`define LDPC_CSR_LDPC_ENC_CODEWRD_VLD_BYTE_OFFSET 13'h03e0
`define LDPC_CSR_LDPC_DEC_SEL_FRMC_SEL_Q0_FRMC_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_SEL_FRMC_SEL_Q0_FRMC_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_SEL_FRMC_SEL_Q0_FRMC_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_SEL_FRMC_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_SEL_FRMC_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_SEL_FRMC_BYTE_OFFSET 13'h03e4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_0_ERR_INTRO_Q0_0_0_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_0_ERR_INTRO_Q0_0_0_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_0_ERR_INTRO_Q0_0_0_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_0_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_0_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_0_BYTE_OFFSET 13'h03e8
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_1_ERR_INTRO_Q0_0_1_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_1_ERR_INTRO_Q0_0_1_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_1_ERR_INTRO_Q0_0_1_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_1_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_1_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_1_BYTE_OFFSET 13'h03ec
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_2_ERR_INTRO_Q0_0_2_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_2_ERR_INTRO_Q0_0_2_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_2_ERR_INTRO_Q0_0_2_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_2_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_2_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_2_BYTE_OFFSET 13'h03f0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_3_ERR_INTRO_Q0_0_3_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_3_ERR_INTRO_Q0_0_3_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_3_ERR_INTRO_Q0_0_3_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_3_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_3_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_3_BYTE_OFFSET 13'h03f4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_4_ERR_INTRO_Q0_0_4_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_4_ERR_INTRO_Q0_0_4_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_4_ERR_INTRO_Q0_0_4_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_4_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_4_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_4_BYTE_OFFSET 13'h03f8
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_5_ERR_INTRO_Q0_0_5_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_5_ERR_INTRO_Q0_0_5_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_5_ERR_INTRO_Q0_0_5_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_5_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_5_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_5_BYTE_OFFSET 13'h03fc
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_6_ERR_INTRO_Q0_0_6_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_6_ERR_INTRO_Q0_0_6_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_6_ERR_INTRO_Q0_0_6_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_6_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_6_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_6_BYTE_OFFSET 13'h0400
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_7_ERR_INTRO_Q0_0_7_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_7_ERR_INTRO_Q0_0_7_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_7_ERR_INTRO_Q0_0_7_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_7_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_7_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_7_BYTE_OFFSET 13'h0404
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_8_ERR_INTRO_Q0_0_8_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_8_ERR_INTRO_Q0_0_8_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_8_ERR_INTRO_Q0_0_8_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_8_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_8_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_8_BYTE_OFFSET 13'h0408
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_9_ERR_INTRO_Q0_0_9_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_9_ERR_INTRO_Q0_0_9_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_9_ERR_INTRO_Q0_0_9_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_9_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_9_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_9_BYTE_OFFSET 13'h040c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_10_ERR_INTRO_Q0_0_10_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_10_ERR_INTRO_Q0_0_10_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_10_ERR_INTRO_Q0_0_10_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_10_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_10_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_10_BYTE_OFFSET 13'h0410
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_11_ERR_INTRO_Q0_0_11_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_11_ERR_INTRO_Q0_0_11_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_11_ERR_INTRO_Q0_0_11_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_11_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_11_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_11_BYTE_OFFSET 13'h0414
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_12_ERR_INTRO_Q0_0_12_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_12_ERR_INTRO_Q0_0_12_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_12_ERR_INTRO_Q0_0_12_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_12_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_12_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_12_BYTE_OFFSET 13'h0418
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_13_ERR_INTRO_Q0_0_13_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_13_ERR_INTRO_Q0_0_13_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_13_ERR_INTRO_Q0_0_13_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_13_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_13_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_13_BYTE_OFFSET 13'h041c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_14_ERR_INTRO_Q0_0_14_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_14_ERR_INTRO_Q0_0_14_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_14_ERR_INTRO_Q0_0_14_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_14_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_14_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_14_BYTE_OFFSET 13'h0420
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_15_ERR_INTRO_Q0_0_15_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_15_ERR_INTRO_Q0_0_15_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_15_ERR_INTRO_Q0_0_15_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_15_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_15_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_15_BYTE_OFFSET 13'h0424
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_16_ERR_INTRO_Q0_0_16_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_16_ERR_INTRO_Q0_0_16_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_16_ERR_INTRO_Q0_0_16_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_16_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_16_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_16_BYTE_OFFSET 13'h0428
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_17_ERR_INTRO_Q0_0_17_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_17_ERR_INTRO_Q0_0_17_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_17_ERR_INTRO_Q0_0_17_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_17_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_17_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_17_BYTE_OFFSET 13'h042c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_18_ERR_INTRO_Q0_0_18_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_18_ERR_INTRO_Q0_0_18_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_18_ERR_INTRO_Q0_0_18_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_18_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_18_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_18_BYTE_OFFSET 13'h0430
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_19_ERR_INTRO_Q0_0_19_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_19_ERR_INTRO_Q0_0_19_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_19_ERR_INTRO_Q0_0_19_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_19_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_19_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_19_BYTE_OFFSET 13'h0434
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_20_ERR_INTRO_Q0_0_20_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_20_ERR_INTRO_Q0_0_20_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_20_ERR_INTRO_Q0_0_20_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_20_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_20_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_20_BYTE_OFFSET 13'h0438
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_21_ERR_INTRO_Q0_0_21_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_21_ERR_INTRO_Q0_0_21_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_21_ERR_INTRO_Q0_0_21_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_21_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_21_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_21_BYTE_OFFSET 13'h043c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_22_ERR_INTRO_Q0_0_22_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_22_ERR_INTRO_Q0_0_22_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_22_ERR_INTRO_Q0_0_22_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_22_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_22_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_22_BYTE_OFFSET 13'h0440
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_23_ERR_INTRO_Q0_0_23_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_23_ERR_INTRO_Q0_0_23_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_23_ERR_INTRO_Q0_0_23_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_23_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_23_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_23_BYTE_OFFSET 13'h0444
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_24_ERR_INTRO_Q0_0_24_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_24_ERR_INTRO_Q0_0_24_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_24_ERR_INTRO_Q0_0_24_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_24_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_24_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_24_BYTE_OFFSET 13'h0448
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_25_ERR_INTRO_Q0_0_25_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_25_ERR_INTRO_Q0_0_25_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_25_ERR_INTRO_Q0_0_25_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_25_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_25_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_25_BYTE_OFFSET 13'h044c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_26_ERR_INTRO_Q0_0_26_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_26_ERR_INTRO_Q0_0_26_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_26_ERR_INTRO_Q0_0_26_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_26_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_26_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_26_BYTE_OFFSET 13'h0450
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_27_ERR_INTRO_Q0_0_27_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_27_ERR_INTRO_Q0_0_27_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_27_ERR_INTRO_Q0_0_27_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_27_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_27_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_27_BYTE_OFFSET 13'h0454
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_28_ERR_INTRO_Q0_0_28_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_28_ERR_INTRO_Q0_0_28_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_28_ERR_INTRO_Q0_0_28_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_28_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_28_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_28_BYTE_OFFSET 13'h0458
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_29_ERR_INTRO_Q0_0_29_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_29_ERR_INTRO_Q0_0_29_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_29_ERR_INTRO_Q0_0_29_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_29_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_29_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_29_BYTE_OFFSET 13'h045c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_30_ERR_INTRO_Q0_0_30_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_30_ERR_INTRO_Q0_0_30_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_30_ERR_INTRO_Q0_0_30_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_30_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_30_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_30_BYTE_OFFSET 13'h0460
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_31_ERR_INTRO_Q0_0_31_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_31_ERR_INTRO_Q0_0_31_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_31_ERR_INTRO_Q0_0_31_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_31_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_31_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_31_BYTE_OFFSET 13'h0464
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_32_ERR_INTRO_Q0_0_32_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_32_ERR_INTRO_Q0_0_32_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_32_ERR_INTRO_Q0_0_32_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_32_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_32_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_32_BYTE_OFFSET 13'h0468
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_33_ERR_INTRO_Q0_0_33_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_33_ERR_INTRO_Q0_0_33_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_33_ERR_INTRO_Q0_0_33_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_33_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_33_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_33_BYTE_OFFSET 13'h046c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_34_ERR_INTRO_Q0_0_34_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_34_ERR_INTRO_Q0_0_34_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_34_ERR_INTRO_Q0_0_34_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_34_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_34_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_34_BYTE_OFFSET 13'h0470
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_35_ERR_INTRO_Q0_0_35_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_35_ERR_INTRO_Q0_0_35_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_35_ERR_INTRO_Q0_0_35_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_35_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_35_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_35_BYTE_OFFSET 13'h0474
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_36_ERR_INTRO_Q0_0_36_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_36_ERR_INTRO_Q0_0_36_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_36_ERR_INTRO_Q0_0_36_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_36_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_36_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_36_BYTE_OFFSET 13'h0478
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_37_ERR_INTRO_Q0_0_37_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_37_ERR_INTRO_Q0_0_37_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_37_ERR_INTRO_Q0_0_37_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_37_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_37_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_37_BYTE_OFFSET 13'h047c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_38_ERR_INTRO_Q0_0_38_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_38_ERR_INTRO_Q0_0_38_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_38_ERR_INTRO_Q0_0_38_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_38_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_38_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_38_BYTE_OFFSET 13'h0480
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_39_ERR_INTRO_Q0_0_39_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_39_ERR_INTRO_Q0_0_39_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_39_ERR_INTRO_Q0_0_39_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_39_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_39_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_39_BYTE_OFFSET 13'h0484
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_40_ERR_INTRO_Q0_0_40_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_40_ERR_INTRO_Q0_0_40_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_40_ERR_INTRO_Q0_0_40_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_40_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_40_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_40_BYTE_OFFSET 13'h0488
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_41_ERR_INTRO_Q0_0_41_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_41_ERR_INTRO_Q0_0_41_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_41_ERR_INTRO_Q0_0_41_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_41_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_41_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_41_BYTE_OFFSET 13'h048c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_42_ERR_INTRO_Q0_0_42_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_42_ERR_INTRO_Q0_0_42_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_42_ERR_INTRO_Q0_0_42_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_42_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_42_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_42_BYTE_OFFSET 13'h0490
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_43_ERR_INTRO_Q0_0_43_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_43_ERR_INTRO_Q0_0_43_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_43_ERR_INTRO_Q0_0_43_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_43_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_43_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_43_BYTE_OFFSET 13'h0494
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_44_ERR_INTRO_Q0_0_44_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_44_ERR_INTRO_Q0_0_44_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_44_ERR_INTRO_Q0_0_44_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_44_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_44_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_44_BYTE_OFFSET 13'h0498
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_45_ERR_INTRO_Q0_0_45_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_45_ERR_INTRO_Q0_0_45_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_45_ERR_INTRO_Q0_0_45_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_45_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_45_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_45_BYTE_OFFSET 13'h049c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_46_ERR_INTRO_Q0_0_46_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_46_ERR_INTRO_Q0_0_46_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_46_ERR_INTRO_Q0_0_46_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_46_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_46_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_46_BYTE_OFFSET 13'h04a0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_47_ERR_INTRO_Q0_0_47_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_47_ERR_INTRO_Q0_0_47_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_47_ERR_INTRO_Q0_0_47_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_47_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_47_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_47_BYTE_OFFSET 13'h04a4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_48_ERR_INTRO_Q0_0_48_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_48_ERR_INTRO_Q0_0_48_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_48_ERR_INTRO_Q0_0_48_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_48_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_48_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_48_BYTE_OFFSET 13'h04a8
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_49_ERR_INTRO_Q0_0_49_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_49_ERR_INTRO_Q0_0_49_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_49_ERR_INTRO_Q0_0_49_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_49_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_49_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_49_BYTE_OFFSET 13'h04ac
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_50_ERR_INTRO_Q0_0_50_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_50_ERR_INTRO_Q0_0_50_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_50_ERR_INTRO_Q0_0_50_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_50_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_50_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_50_BYTE_OFFSET 13'h04b0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_51_ERR_INTRO_Q0_0_51_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_51_ERR_INTRO_Q0_0_51_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_51_ERR_INTRO_Q0_0_51_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_51_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_51_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_51_BYTE_OFFSET 13'h04b4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_52_ERR_INTRO_Q0_0_52_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_52_ERR_INTRO_Q0_0_52_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_52_ERR_INTRO_Q0_0_52_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_52_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_52_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_52_BYTE_OFFSET 13'h04b8
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_53_ERR_INTRO_Q0_0_53_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_53_ERR_INTRO_Q0_0_53_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_53_ERR_INTRO_Q0_0_53_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_53_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_53_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_53_BYTE_OFFSET 13'h04bc
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_54_ERR_INTRO_Q0_0_54_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_54_ERR_INTRO_Q0_0_54_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_54_ERR_INTRO_Q0_0_54_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_54_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_54_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_54_BYTE_OFFSET 13'h04c0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_55_ERR_INTRO_Q0_0_55_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_55_ERR_INTRO_Q0_0_55_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_55_ERR_INTRO_Q0_0_55_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_55_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_55_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_55_BYTE_OFFSET 13'h04c4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_56_ERR_INTRO_Q0_0_56_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_56_ERR_INTRO_Q0_0_56_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_56_ERR_INTRO_Q0_0_56_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_56_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_56_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_56_BYTE_OFFSET 13'h04c8
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_57_ERR_INTRO_Q0_0_57_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_57_ERR_INTRO_Q0_0_57_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_57_ERR_INTRO_Q0_0_57_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_57_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_57_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_57_BYTE_OFFSET 13'h04cc
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_58_ERR_INTRO_Q0_0_58_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_58_ERR_INTRO_Q0_0_58_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_58_ERR_INTRO_Q0_0_58_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_58_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_58_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_58_BYTE_OFFSET 13'h04d0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_59_ERR_INTRO_Q0_0_59_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_59_ERR_INTRO_Q0_0_59_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_59_ERR_INTRO_Q0_0_59_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_59_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_59_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_59_BYTE_OFFSET 13'h04d4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_60_ERR_INTRO_Q0_0_60_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_60_ERR_INTRO_Q0_0_60_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_60_ERR_INTRO_Q0_0_60_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_60_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_60_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_60_BYTE_OFFSET 13'h04d8
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_61_ERR_INTRO_Q0_0_61_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_61_ERR_INTRO_Q0_0_61_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_61_ERR_INTRO_Q0_0_61_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_61_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_61_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_61_BYTE_OFFSET 13'h04dc
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_62_ERR_INTRO_Q0_0_62_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_62_ERR_INTRO_Q0_0_62_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_62_ERR_INTRO_Q0_0_62_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_62_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_62_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_62_BYTE_OFFSET 13'h04e0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_63_ERR_INTRO_Q0_0_63_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_63_ERR_INTRO_Q0_0_63_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_63_ERR_INTRO_Q0_0_63_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_63_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_63_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_63_BYTE_OFFSET 13'h04e4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_64_ERR_INTRO_Q0_0_64_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_64_ERR_INTRO_Q0_0_64_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_64_ERR_INTRO_Q0_0_64_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_64_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_64_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_64_BYTE_OFFSET 13'h04e8
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_65_ERR_INTRO_Q0_0_65_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_65_ERR_INTRO_Q0_0_65_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_65_ERR_INTRO_Q0_0_65_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_65_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_65_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_65_BYTE_OFFSET 13'h04ec
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_66_ERR_INTRO_Q0_0_66_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_66_ERR_INTRO_Q0_0_66_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_66_ERR_INTRO_Q0_0_66_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_66_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_66_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_66_BYTE_OFFSET 13'h04f0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_67_ERR_INTRO_Q0_0_67_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_67_ERR_INTRO_Q0_0_67_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_67_ERR_INTRO_Q0_0_67_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_67_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_67_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_67_BYTE_OFFSET 13'h04f4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_68_ERR_INTRO_Q0_0_68_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_68_ERR_INTRO_Q0_0_68_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_68_ERR_INTRO_Q0_0_68_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_68_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_68_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_68_BYTE_OFFSET 13'h04f8
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_69_ERR_INTRO_Q0_0_69_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_69_ERR_INTRO_Q0_0_69_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_69_ERR_INTRO_Q0_0_69_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_69_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_69_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_69_BYTE_OFFSET 13'h04fc
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_70_ERR_INTRO_Q0_0_70_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_70_ERR_INTRO_Q0_0_70_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_70_ERR_INTRO_Q0_0_70_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_70_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_70_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_70_BYTE_OFFSET 13'h0500
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_71_ERR_INTRO_Q0_0_71_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_71_ERR_INTRO_Q0_0_71_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_71_ERR_INTRO_Q0_0_71_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_71_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_71_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_71_BYTE_OFFSET 13'h0504
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_72_ERR_INTRO_Q0_0_72_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_72_ERR_INTRO_Q0_0_72_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_72_ERR_INTRO_Q0_0_72_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_72_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_72_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_72_BYTE_OFFSET 13'h0508
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_73_ERR_INTRO_Q0_0_73_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_73_ERR_INTRO_Q0_0_73_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_73_ERR_INTRO_Q0_0_73_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_73_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_73_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_73_BYTE_OFFSET 13'h050c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_74_ERR_INTRO_Q0_0_74_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_74_ERR_INTRO_Q0_0_74_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_74_ERR_INTRO_Q0_0_74_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_74_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_74_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_74_BYTE_OFFSET 13'h0510
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_75_ERR_INTRO_Q0_0_75_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_75_ERR_INTRO_Q0_0_75_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_75_ERR_INTRO_Q0_0_75_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_75_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_75_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_75_BYTE_OFFSET 13'h0514
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_76_ERR_INTRO_Q0_0_76_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_76_ERR_INTRO_Q0_0_76_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_76_ERR_INTRO_Q0_0_76_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_76_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_76_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_76_BYTE_OFFSET 13'h0518
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_77_ERR_INTRO_Q0_0_77_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_77_ERR_INTRO_Q0_0_77_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_77_ERR_INTRO_Q0_0_77_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_77_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_77_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_77_BYTE_OFFSET 13'h051c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_78_ERR_INTRO_Q0_0_78_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_78_ERR_INTRO_Q0_0_78_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_78_ERR_INTRO_Q0_0_78_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_78_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_78_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_78_BYTE_OFFSET 13'h0520
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_79_ERR_INTRO_Q0_0_79_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_79_ERR_INTRO_Q0_0_79_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_79_ERR_INTRO_Q0_0_79_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_79_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_79_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_79_BYTE_OFFSET 13'h0524
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_80_ERR_INTRO_Q0_0_80_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_80_ERR_INTRO_Q0_0_80_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_80_ERR_INTRO_Q0_0_80_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_80_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_80_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_80_BYTE_OFFSET 13'h0528
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_81_ERR_INTRO_Q0_0_81_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_81_ERR_INTRO_Q0_0_81_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_81_ERR_INTRO_Q0_0_81_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_81_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_81_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_81_BYTE_OFFSET 13'h052c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_82_ERR_INTRO_Q0_0_82_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_82_ERR_INTRO_Q0_0_82_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_82_ERR_INTRO_Q0_0_82_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_82_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_82_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_82_BYTE_OFFSET 13'h0530
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_83_ERR_INTRO_Q0_0_83_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_83_ERR_INTRO_Q0_0_83_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_83_ERR_INTRO_Q0_0_83_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_83_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_83_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_83_BYTE_OFFSET 13'h0534
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_84_ERR_INTRO_Q0_0_84_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_84_ERR_INTRO_Q0_0_84_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_84_ERR_INTRO_Q0_0_84_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_84_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_84_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_84_BYTE_OFFSET 13'h0538
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_85_ERR_INTRO_Q0_0_85_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_85_ERR_INTRO_Q0_0_85_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_85_ERR_INTRO_Q0_0_85_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_85_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_85_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_85_BYTE_OFFSET 13'h053c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_86_ERR_INTRO_Q0_0_86_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_86_ERR_INTRO_Q0_0_86_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_86_ERR_INTRO_Q0_0_86_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_86_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_86_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_86_BYTE_OFFSET 13'h0540
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_87_ERR_INTRO_Q0_0_87_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_87_ERR_INTRO_Q0_0_87_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_87_ERR_INTRO_Q0_0_87_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_87_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_87_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_87_BYTE_OFFSET 13'h0544
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_88_ERR_INTRO_Q0_0_88_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_88_ERR_INTRO_Q0_0_88_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_88_ERR_INTRO_Q0_0_88_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_88_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_88_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_88_BYTE_OFFSET 13'h0548
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_89_ERR_INTRO_Q0_0_89_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_89_ERR_INTRO_Q0_0_89_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_89_ERR_INTRO_Q0_0_89_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_89_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_89_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_89_BYTE_OFFSET 13'h054c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_90_ERR_INTRO_Q0_0_90_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_90_ERR_INTRO_Q0_0_90_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_90_ERR_INTRO_Q0_0_90_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_90_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_90_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_90_BYTE_OFFSET 13'h0550
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_91_ERR_INTRO_Q0_0_91_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_91_ERR_INTRO_Q0_0_91_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_91_ERR_INTRO_Q0_0_91_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_91_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_91_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_91_BYTE_OFFSET 13'h0554
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_92_ERR_INTRO_Q0_0_92_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_92_ERR_INTRO_Q0_0_92_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_92_ERR_INTRO_Q0_0_92_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_92_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_92_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_92_BYTE_OFFSET 13'h0558
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_93_ERR_INTRO_Q0_0_93_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_93_ERR_INTRO_Q0_0_93_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_93_ERR_INTRO_Q0_0_93_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_93_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_93_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_93_BYTE_OFFSET 13'h055c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_94_ERR_INTRO_Q0_0_94_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_94_ERR_INTRO_Q0_0_94_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_94_ERR_INTRO_Q0_0_94_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_94_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_94_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_94_BYTE_OFFSET 13'h0560
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_95_ERR_INTRO_Q0_0_95_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_95_ERR_INTRO_Q0_0_95_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_95_ERR_INTRO_Q0_0_95_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_95_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_95_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_95_BYTE_OFFSET 13'h0564
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_96_ERR_INTRO_Q0_0_96_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_96_ERR_INTRO_Q0_0_96_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_96_ERR_INTRO_Q0_0_96_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_96_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_96_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_96_BYTE_OFFSET 13'h0568
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_97_ERR_INTRO_Q0_0_97_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_97_ERR_INTRO_Q0_0_97_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_97_ERR_INTRO_Q0_0_97_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_97_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_97_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_97_BYTE_OFFSET 13'h056c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_98_ERR_INTRO_Q0_0_98_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_98_ERR_INTRO_Q0_0_98_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_98_ERR_INTRO_Q0_0_98_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_98_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_98_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_98_BYTE_OFFSET 13'h0570
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_99_ERR_INTRO_Q0_0_99_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_99_ERR_INTRO_Q0_0_99_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_99_ERR_INTRO_Q0_0_99_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_99_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_99_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_99_BYTE_OFFSET 13'h0574
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_100_ERR_INTRO_Q0_0_100_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_100_ERR_INTRO_Q0_0_100_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_100_ERR_INTRO_Q0_0_100_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_100_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_100_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_100_BYTE_OFFSET 13'h0578
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_101_ERR_INTRO_Q0_0_101_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_101_ERR_INTRO_Q0_0_101_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_101_ERR_INTRO_Q0_0_101_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_101_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_101_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_101_BYTE_OFFSET 13'h057c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_102_ERR_INTRO_Q0_0_102_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_102_ERR_INTRO_Q0_0_102_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_102_ERR_INTRO_Q0_0_102_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_102_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_102_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_102_BYTE_OFFSET 13'h0580
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_103_ERR_INTRO_Q0_0_103_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_103_ERR_INTRO_Q0_0_103_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_103_ERR_INTRO_Q0_0_103_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_103_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_103_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_103_BYTE_OFFSET 13'h0584
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_104_ERR_INTRO_Q0_0_104_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_104_ERR_INTRO_Q0_0_104_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_104_ERR_INTRO_Q0_0_104_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_104_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_104_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_104_BYTE_OFFSET 13'h0588
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_105_ERR_INTRO_Q0_0_105_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_105_ERR_INTRO_Q0_0_105_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_105_ERR_INTRO_Q0_0_105_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_105_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_105_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_105_BYTE_OFFSET 13'h058c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_106_ERR_INTRO_Q0_0_106_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_106_ERR_INTRO_Q0_0_106_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_106_ERR_INTRO_Q0_0_106_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_106_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_106_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_106_BYTE_OFFSET 13'h0590
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_107_ERR_INTRO_Q0_0_107_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_107_ERR_INTRO_Q0_0_107_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_107_ERR_INTRO_Q0_0_107_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_107_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_107_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_107_BYTE_OFFSET 13'h0594
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_108_ERR_INTRO_Q0_0_108_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_108_ERR_INTRO_Q0_0_108_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_108_ERR_INTRO_Q0_0_108_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_108_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_108_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_108_BYTE_OFFSET 13'h0598
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_109_ERR_INTRO_Q0_0_109_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_109_ERR_INTRO_Q0_0_109_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_109_ERR_INTRO_Q0_0_109_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_109_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_109_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_109_BYTE_OFFSET 13'h059c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_110_ERR_INTRO_Q0_0_110_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_110_ERR_INTRO_Q0_0_110_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_110_ERR_INTRO_Q0_0_110_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_110_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_110_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_110_BYTE_OFFSET 13'h05a0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_111_ERR_INTRO_Q0_0_111_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_111_ERR_INTRO_Q0_0_111_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_111_ERR_INTRO_Q0_0_111_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_111_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_111_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_111_BYTE_OFFSET 13'h05a4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_112_ERR_INTRO_Q0_0_112_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_112_ERR_INTRO_Q0_0_112_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_112_ERR_INTRO_Q0_0_112_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_112_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_112_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_112_BYTE_OFFSET 13'h05a8
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_113_ERR_INTRO_Q0_0_113_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_113_ERR_INTRO_Q0_0_113_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_113_ERR_INTRO_Q0_0_113_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_113_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_113_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_113_BYTE_OFFSET 13'h05ac
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_114_ERR_INTRO_Q0_0_114_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_114_ERR_INTRO_Q0_0_114_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_114_ERR_INTRO_Q0_0_114_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_114_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_114_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_114_BYTE_OFFSET 13'h05b0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_115_ERR_INTRO_Q0_0_115_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_115_ERR_INTRO_Q0_0_115_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_115_ERR_INTRO_Q0_0_115_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_115_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_115_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_115_BYTE_OFFSET 13'h05b4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_116_ERR_INTRO_Q0_0_116_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_116_ERR_INTRO_Q0_0_116_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_116_ERR_INTRO_Q0_0_116_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_116_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_116_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_116_BYTE_OFFSET 13'h05b8
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_117_ERR_INTRO_Q0_0_117_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_117_ERR_INTRO_Q0_0_117_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_117_ERR_INTRO_Q0_0_117_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_117_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_117_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_117_BYTE_OFFSET 13'h05bc
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_118_ERR_INTRO_Q0_0_118_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_118_ERR_INTRO_Q0_0_118_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_118_ERR_INTRO_Q0_0_118_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_118_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_118_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_118_BYTE_OFFSET 13'h05c0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_119_ERR_INTRO_Q0_0_119_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_119_ERR_INTRO_Q0_0_119_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_119_ERR_INTRO_Q0_0_119_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_119_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_119_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_119_BYTE_OFFSET 13'h05c4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_120_ERR_INTRO_Q0_0_120_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_120_ERR_INTRO_Q0_0_120_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_120_ERR_INTRO_Q0_0_120_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_120_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_120_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_120_BYTE_OFFSET 13'h05c8
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_121_ERR_INTRO_Q0_0_121_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_121_ERR_INTRO_Q0_0_121_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_121_ERR_INTRO_Q0_0_121_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_121_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_121_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_121_BYTE_OFFSET 13'h05cc
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_122_ERR_INTRO_Q0_0_122_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_122_ERR_INTRO_Q0_0_122_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_122_ERR_INTRO_Q0_0_122_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_122_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_122_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_122_BYTE_OFFSET 13'h05d0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_123_ERR_INTRO_Q0_0_123_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_123_ERR_INTRO_Q0_0_123_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_123_ERR_INTRO_Q0_0_123_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_123_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_123_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_123_BYTE_OFFSET 13'h05d4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_124_ERR_INTRO_Q0_0_124_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_124_ERR_INTRO_Q0_0_124_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_124_ERR_INTRO_Q0_0_124_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_124_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_124_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_124_BYTE_OFFSET 13'h05d8
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_125_ERR_INTRO_Q0_0_125_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_125_ERR_INTRO_Q0_0_125_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_125_ERR_INTRO_Q0_0_125_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_125_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_125_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_125_BYTE_OFFSET 13'h05dc
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_126_ERR_INTRO_Q0_0_126_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_126_ERR_INTRO_Q0_0_126_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_126_ERR_INTRO_Q0_0_126_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_126_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_126_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_126_BYTE_OFFSET 13'h05e0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_127_ERR_INTRO_Q0_0_127_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_127_ERR_INTRO_Q0_0_127_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_127_ERR_INTRO_Q0_0_127_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_127_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_127_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_127_BYTE_OFFSET 13'h05e4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_128_ERR_INTRO_Q0_0_128_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_128_ERR_INTRO_Q0_0_128_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_128_ERR_INTRO_Q0_0_128_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_128_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_128_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_128_BYTE_OFFSET 13'h05e8
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_129_ERR_INTRO_Q0_0_129_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_129_ERR_INTRO_Q0_0_129_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_129_ERR_INTRO_Q0_0_129_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_129_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_129_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_129_BYTE_OFFSET 13'h05ec
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_130_ERR_INTRO_Q0_0_130_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_130_ERR_INTRO_Q0_0_130_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_130_ERR_INTRO_Q0_0_130_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_130_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_130_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_130_BYTE_OFFSET 13'h05f0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_131_ERR_INTRO_Q0_0_131_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_131_ERR_INTRO_Q0_0_131_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_131_ERR_INTRO_Q0_0_131_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_131_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_131_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_131_BYTE_OFFSET 13'h05f4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_132_ERR_INTRO_Q0_0_132_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_132_ERR_INTRO_Q0_0_132_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_132_ERR_INTRO_Q0_0_132_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_132_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_132_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_132_BYTE_OFFSET 13'h05f8
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_133_ERR_INTRO_Q0_0_133_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_133_ERR_INTRO_Q0_0_133_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_133_ERR_INTRO_Q0_0_133_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_133_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_133_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_133_BYTE_OFFSET 13'h05fc
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_134_ERR_INTRO_Q0_0_134_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_134_ERR_INTRO_Q0_0_134_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_134_ERR_INTRO_Q0_0_134_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_134_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_134_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_134_BYTE_OFFSET 13'h0600
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_135_ERR_INTRO_Q0_0_135_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_135_ERR_INTRO_Q0_0_135_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_135_ERR_INTRO_Q0_0_135_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_135_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_135_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_135_BYTE_OFFSET 13'h0604
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_136_ERR_INTRO_Q0_0_136_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_136_ERR_INTRO_Q0_0_136_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_136_ERR_INTRO_Q0_0_136_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_136_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_136_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_136_BYTE_OFFSET 13'h0608
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_137_ERR_INTRO_Q0_0_137_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_137_ERR_INTRO_Q0_0_137_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_137_ERR_INTRO_Q0_0_137_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_137_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_137_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_137_BYTE_OFFSET 13'h060c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_138_ERR_INTRO_Q0_0_138_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_138_ERR_INTRO_Q0_0_138_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_138_ERR_INTRO_Q0_0_138_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_138_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_138_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_138_BYTE_OFFSET 13'h0610
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_139_ERR_INTRO_Q0_0_139_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_139_ERR_INTRO_Q0_0_139_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_139_ERR_INTRO_Q0_0_139_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_139_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_139_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_139_BYTE_OFFSET 13'h0614
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_140_ERR_INTRO_Q0_0_140_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_140_ERR_INTRO_Q0_0_140_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_140_ERR_INTRO_Q0_0_140_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_140_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_140_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_140_BYTE_OFFSET 13'h0618
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_141_ERR_INTRO_Q0_0_141_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_141_ERR_INTRO_Q0_0_141_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_141_ERR_INTRO_Q0_0_141_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_141_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_141_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_141_BYTE_OFFSET 13'h061c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_142_ERR_INTRO_Q0_0_142_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_142_ERR_INTRO_Q0_0_142_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_142_ERR_INTRO_Q0_0_142_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_142_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_142_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_142_BYTE_OFFSET 13'h0620
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_143_ERR_INTRO_Q0_0_143_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_143_ERR_INTRO_Q0_0_143_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_143_ERR_INTRO_Q0_0_143_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_143_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_143_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_143_BYTE_OFFSET 13'h0624
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_144_ERR_INTRO_Q0_0_144_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_144_ERR_INTRO_Q0_0_144_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_144_ERR_INTRO_Q0_0_144_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_144_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_144_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_144_BYTE_OFFSET 13'h0628
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_145_ERR_INTRO_Q0_0_145_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_145_ERR_INTRO_Q0_0_145_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_145_ERR_INTRO_Q0_0_145_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_145_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_145_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_145_BYTE_OFFSET 13'h062c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_146_ERR_INTRO_Q0_0_146_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_146_ERR_INTRO_Q0_0_146_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_146_ERR_INTRO_Q0_0_146_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_146_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_146_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_146_BYTE_OFFSET 13'h0630
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_147_ERR_INTRO_Q0_0_147_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_147_ERR_INTRO_Q0_0_147_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_147_ERR_INTRO_Q0_0_147_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_147_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_147_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_147_BYTE_OFFSET 13'h0634
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_148_ERR_INTRO_Q0_0_148_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_148_ERR_INTRO_Q0_0_148_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_148_ERR_INTRO_Q0_0_148_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_148_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_148_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_148_BYTE_OFFSET 13'h0638
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_149_ERR_INTRO_Q0_0_149_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_149_ERR_INTRO_Q0_0_149_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_149_ERR_INTRO_Q0_0_149_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_149_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_149_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_149_BYTE_OFFSET 13'h063c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_150_ERR_INTRO_Q0_0_150_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_150_ERR_INTRO_Q0_0_150_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_150_ERR_INTRO_Q0_0_150_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_150_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_150_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_150_BYTE_OFFSET 13'h0640
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_151_ERR_INTRO_Q0_0_151_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_151_ERR_INTRO_Q0_0_151_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_151_ERR_INTRO_Q0_0_151_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_151_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_151_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_151_BYTE_OFFSET 13'h0644
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_152_ERR_INTRO_Q0_0_152_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_152_ERR_INTRO_Q0_0_152_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_152_ERR_INTRO_Q0_0_152_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_152_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_152_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_152_BYTE_OFFSET 13'h0648
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_153_ERR_INTRO_Q0_0_153_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_153_ERR_INTRO_Q0_0_153_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_153_ERR_INTRO_Q0_0_153_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_153_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_153_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_153_BYTE_OFFSET 13'h064c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_154_ERR_INTRO_Q0_0_154_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_154_ERR_INTRO_Q0_0_154_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_154_ERR_INTRO_Q0_0_154_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_154_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_154_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_154_BYTE_OFFSET 13'h0650
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_155_ERR_INTRO_Q0_0_155_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_155_ERR_INTRO_Q0_0_155_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_155_ERR_INTRO_Q0_0_155_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_155_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_155_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_155_BYTE_OFFSET 13'h0654
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_156_ERR_INTRO_Q0_0_156_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_156_ERR_INTRO_Q0_0_156_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_156_ERR_INTRO_Q0_0_156_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_156_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_156_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_156_BYTE_OFFSET 13'h0658
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_157_ERR_INTRO_Q0_0_157_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_157_ERR_INTRO_Q0_0_157_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_157_ERR_INTRO_Q0_0_157_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_157_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_157_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_157_BYTE_OFFSET 13'h065c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_158_ERR_INTRO_Q0_0_158_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_158_ERR_INTRO_Q0_0_158_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_158_ERR_INTRO_Q0_0_158_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_158_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_158_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_158_BYTE_OFFSET 13'h0660
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_159_ERR_INTRO_Q0_0_159_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_159_ERR_INTRO_Q0_0_159_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_159_ERR_INTRO_Q0_0_159_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_159_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_159_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_159_BYTE_OFFSET 13'h0664
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_160_ERR_INTRO_Q0_0_160_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_160_ERR_INTRO_Q0_0_160_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_160_ERR_INTRO_Q0_0_160_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_160_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_160_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_160_BYTE_OFFSET 13'h0668
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_161_ERR_INTRO_Q0_0_161_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_161_ERR_INTRO_Q0_0_161_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_161_ERR_INTRO_Q0_0_161_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_161_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_161_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_161_BYTE_OFFSET 13'h066c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_162_ERR_INTRO_Q0_0_162_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_162_ERR_INTRO_Q0_0_162_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_162_ERR_INTRO_Q0_0_162_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_162_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_162_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_162_BYTE_OFFSET 13'h0670
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_163_ERR_INTRO_Q0_0_163_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_163_ERR_INTRO_Q0_0_163_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_163_ERR_INTRO_Q0_0_163_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_163_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_163_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_163_BYTE_OFFSET 13'h0674
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_164_ERR_INTRO_Q0_0_164_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_164_ERR_INTRO_Q0_0_164_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_164_ERR_INTRO_Q0_0_164_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_164_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_164_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_164_BYTE_OFFSET 13'h0678
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_165_ERR_INTRO_Q0_0_165_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_165_ERR_INTRO_Q0_0_165_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_165_ERR_INTRO_Q0_0_165_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_165_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_165_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_165_BYTE_OFFSET 13'h067c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_166_ERR_INTRO_Q0_0_166_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_166_ERR_INTRO_Q0_0_166_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_166_ERR_INTRO_Q0_0_166_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_166_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_166_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_166_BYTE_OFFSET 13'h0680
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_167_ERR_INTRO_Q0_0_167_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_167_ERR_INTRO_Q0_0_167_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_167_ERR_INTRO_Q0_0_167_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_167_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_167_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_167_BYTE_OFFSET 13'h0684
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_168_ERR_INTRO_Q0_0_168_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_168_ERR_INTRO_Q0_0_168_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_168_ERR_INTRO_Q0_0_168_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_168_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_168_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_168_BYTE_OFFSET 13'h0688
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_169_ERR_INTRO_Q0_0_169_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_169_ERR_INTRO_Q0_0_169_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_169_ERR_INTRO_Q0_0_169_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_169_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_169_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_169_BYTE_OFFSET 13'h068c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_170_ERR_INTRO_Q0_0_170_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_170_ERR_INTRO_Q0_0_170_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_170_ERR_INTRO_Q0_0_170_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_170_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_170_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_170_BYTE_OFFSET 13'h0690
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_171_ERR_INTRO_Q0_0_171_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_171_ERR_INTRO_Q0_0_171_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_171_ERR_INTRO_Q0_0_171_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_171_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_171_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_171_BYTE_OFFSET 13'h0694
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_172_ERR_INTRO_Q0_0_172_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_172_ERR_INTRO_Q0_0_172_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_172_ERR_INTRO_Q0_0_172_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_172_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_172_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_172_BYTE_OFFSET 13'h0698
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_173_ERR_INTRO_Q0_0_173_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_173_ERR_INTRO_Q0_0_173_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_173_ERR_INTRO_Q0_0_173_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_173_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_173_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_173_BYTE_OFFSET 13'h069c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_174_ERR_INTRO_Q0_0_174_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_174_ERR_INTRO_Q0_0_174_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_174_ERR_INTRO_Q0_0_174_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_174_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_174_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_174_BYTE_OFFSET 13'h06a0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_175_ERR_INTRO_Q0_0_175_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_175_ERR_INTRO_Q0_0_175_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_175_ERR_INTRO_Q0_0_175_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_175_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_175_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_175_BYTE_OFFSET 13'h06a4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_176_ERR_INTRO_Q0_0_176_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_176_ERR_INTRO_Q0_0_176_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_176_ERR_INTRO_Q0_0_176_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_176_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_176_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_176_BYTE_OFFSET 13'h06a8
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_177_ERR_INTRO_Q0_0_177_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_177_ERR_INTRO_Q0_0_177_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_177_ERR_INTRO_Q0_0_177_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_177_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_177_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_177_BYTE_OFFSET 13'h06ac
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_178_ERR_INTRO_Q0_0_178_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_178_ERR_INTRO_Q0_0_178_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_178_ERR_INTRO_Q0_0_178_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_178_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_178_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_178_BYTE_OFFSET 13'h06b0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_179_ERR_INTRO_Q0_0_179_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_179_ERR_INTRO_Q0_0_179_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_179_ERR_INTRO_Q0_0_179_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_179_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_179_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_179_BYTE_OFFSET 13'h06b4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_180_ERR_INTRO_Q0_0_180_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_180_ERR_INTRO_Q0_0_180_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_180_ERR_INTRO_Q0_0_180_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_180_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_180_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_180_BYTE_OFFSET 13'h06b8
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_181_ERR_INTRO_Q0_0_181_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_181_ERR_INTRO_Q0_0_181_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_181_ERR_INTRO_Q0_0_181_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_181_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_181_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_181_BYTE_OFFSET 13'h06bc
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_182_ERR_INTRO_Q0_0_182_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_182_ERR_INTRO_Q0_0_182_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_182_ERR_INTRO_Q0_0_182_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_182_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_182_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_182_BYTE_OFFSET 13'h06c0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_183_ERR_INTRO_Q0_0_183_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_183_ERR_INTRO_Q0_0_183_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_183_ERR_INTRO_Q0_0_183_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_183_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_183_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_183_BYTE_OFFSET 13'h06c4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_184_ERR_INTRO_Q0_0_184_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_184_ERR_INTRO_Q0_0_184_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_184_ERR_INTRO_Q0_0_184_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_184_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_184_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_184_BYTE_OFFSET 13'h06c8
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_185_ERR_INTRO_Q0_0_185_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_185_ERR_INTRO_Q0_0_185_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_185_ERR_INTRO_Q0_0_185_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_185_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_185_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_185_BYTE_OFFSET 13'h06cc
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_186_ERR_INTRO_Q0_0_186_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_186_ERR_INTRO_Q0_0_186_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_186_ERR_INTRO_Q0_0_186_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_186_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_186_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_186_BYTE_OFFSET 13'h06d0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_187_ERR_INTRO_Q0_0_187_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_187_ERR_INTRO_Q0_0_187_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_187_ERR_INTRO_Q0_0_187_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_187_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_187_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_187_BYTE_OFFSET 13'h06d4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_188_ERR_INTRO_Q0_0_188_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_188_ERR_INTRO_Q0_0_188_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_188_ERR_INTRO_Q0_0_188_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_188_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_188_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_188_BYTE_OFFSET 13'h06d8
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_189_ERR_INTRO_Q0_0_189_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_189_ERR_INTRO_Q0_0_189_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_189_ERR_INTRO_Q0_0_189_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_189_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_189_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_189_BYTE_OFFSET 13'h06dc
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_190_ERR_INTRO_Q0_0_190_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_190_ERR_INTRO_Q0_0_190_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_190_ERR_INTRO_Q0_0_190_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_190_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_190_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_190_BYTE_OFFSET 13'h06e0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_191_ERR_INTRO_Q0_0_191_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_191_ERR_INTRO_Q0_0_191_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_191_ERR_INTRO_Q0_0_191_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_191_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_191_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_191_BYTE_OFFSET 13'h06e4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_192_ERR_INTRO_Q0_0_192_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_192_ERR_INTRO_Q0_0_192_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_192_ERR_INTRO_Q0_0_192_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_192_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_192_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_192_BYTE_OFFSET 13'h06e8
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_193_ERR_INTRO_Q0_0_193_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_193_ERR_INTRO_Q0_0_193_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_193_ERR_INTRO_Q0_0_193_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_193_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_193_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_193_BYTE_OFFSET 13'h06ec
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_194_ERR_INTRO_Q0_0_194_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_194_ERR_INTRO_Q0_0_194_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_194_ERR_INTRO_Q0_0_194_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_194_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_194_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_194_BYTE_OFFSET 13'h06f0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_195_ERR_INTRO_Q0_0_195_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_195_ERR_INTRO_Q0_0_195_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_195_ERR_INTRO_Q0_0_195_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_195_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_195_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_195_BYTE_OFFSET 13'h06f4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_196_ERR_INTRO_Q0_0_196_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_196_ERR_INTRO_Q0_0_196_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_196_ERR_INTRO_Q0_0_196_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_196_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_196_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_196_BYTE_OFFSET 13'h06f8
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_197_ERR_INTRO_Q0_0_197_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_197_ERR_INTRO_Q0_0_197_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_197_ERR_INTRO_Q0_0_197_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_197_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_197_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_197_BYTE_OFFSET 13'h06fc
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_198_ERR_INTRO_Q0_0_198_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_198_ERR_INTRO_Q0_0_198_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_198_ERR_INTRO_Q0_0_198_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_198_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_198_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_198_BYTE_OFFSET 13'h0700
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_199_ERR_INTRO_Q0_0_199_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_199_ERR_INTRO_Q0_0_199_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_199_ERR_INTRO_Q0_0_199_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_199_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_199_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_199_BYTE_OFFSET 13'h0704
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_200_ERR_INTRO_Q0_0_200_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_200_ERR_INTRO_Q0_0_200_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_200_ERR_INTRO_Q0_0_200_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_200_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_200_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_200_BYTE_OFFSET 13'h0708
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_201_ERR_INTRO_Q0_0_201_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_201_ERR_INTRO_Q0_0_201_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_201_ERR_INTRO_Q0_0_201_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_201_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_201_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_201_BYTE_OFFSET 13'h070c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_202_ERR_INTRO_Q0_0_202_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_202_ERR_INTRO_Q0_0_202_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_202_ERR_INTRO_Q0_0_202_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_202_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_202_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_202_BYTE_OFFSET 13'h0710
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_203_ERR_INTRO_Q0_0_203_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_203_ERR_INTRO_Q0_0_203_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_203_ERR_INTRO_Q0_0_203_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_203_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_203_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_203_BYTE_OFFSET 13'h0714
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_204_ERR_INTRO_Q0_0_204_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_204_ERR_INTRO_Q0_0_204_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_204_ERR_INTRO_Q0_0_204_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_204_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_204_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_204_BYTE_OFFSET 13'h0718
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_205_ERR_INTRO_Q0_0_205_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_205_ERR_INTRO_Q0_0_205_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_205_ERR_INTRO_Q0_0_205_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_205_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_205_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_205_BYTE_OFFSET 13'h071c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_206_ERR_INTRO_Q0_0_206_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_206_ERR_INTRO_Q0_0_206_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_206_ERR_INTRO_Q0_0_206_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_206_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_206_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_206_BYTE_OFFSET 13'h0720
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_207_ERR_INTRO_Q0_0_207_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_207_ERR_INTRO_Q0_0_207_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_207_ERR_INTRO_Q0_0_207_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_207_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_207_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_0_INTRO_207_BYTE_OFFSET 13'h0724
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_0_ERR_INTRO_Q0_1_0_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_0_ERR_INTRO_Q0_1_0_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_0_ERR_INTRO_Q0_1_0_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_0_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_0_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_0_BYTE_OFFSET 13'h0728
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_1_ERR_INTRO_Q0_1_1_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_1_ERR_INTRO_Q0_1_1_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_1_ERR_INTRO_Q0_1_1_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_1_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_1_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_1_BYTE_OFFSET 13'h072c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_2_ERR_INTRO_Q0_1_2_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_2_ERR_INTRO_Q0_1_2_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_2_ERR_INTRO_Q0_1_2_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_2_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_2_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_2_BYTE_OFFSET 13'h0730
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_3_ERR_INTRO_Q0_1_3_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_3_ERR_INTRO_Q0_1_3_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_3_ERR_INTRO_Q0_1_3_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_3_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_3_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_3_BYTE_OFFSET 13'h0734
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_4_ERR_INTRO_Q0_1_4_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_4_ERR_INTRO_Q0_1_4_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_4_ERR_INTRO_Q0_1_4_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_4_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_4_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_4_BYTE_OFFSET 13'h0738
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_5_ERR_INTRO_Q0_1_5_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_5_ERR_INTRO_Q0_1_5_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_5_ERR_INTRO_Q0_1_5_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_5_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_5_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_5_BYTE_OFFSET 13'h073c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_6_ERR_INTRO_Q0_1_6_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_6_ERR_INTRO_Q0_1_6_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_6_ERR_INTRO_Q0_1_6_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_6_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_6_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_6_BYTE_OFFSET 13'h0740
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_7_ERR_INTRO_Q0_1_7_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_7_ERR_INTRO_Q0_1_7_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_7_ERR_INTRO_Q0_1_7_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_7_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_7_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_7_BYTE_OFFSET 13'h0744
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_8_ERR_INTRO_Q0_1_8_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_8_ERR_INTRO_Q0_1_8_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_8_ERR_INTRO_Q0_1_8_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_8_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_8_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_8_BYTE_OFFSET 13'h0748
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_9_ERR_INTRO_Q0_1_9_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_9_ERR_INTRO_Q0_1_9_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_9_ERR_INTRO_Q0_1_9_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_9_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_9_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_9_BYTE_OFFSET 13'h074c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_10_ERR_INTRO_Q0_1_10_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_10_ERR_INTRO_Q0_1_10_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_10_ERR_INTRO_Q0_1_10_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_10_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_10_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_10_BYTE_OFFSET 13'h0750
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_11_ERR_INTRO_Q0_1_11_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_11_ERR_INTRO_Q0_1_11_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_11_ERR_INTRO_Q0_1_11_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_11_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_11_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_11_BYTE_OFFSET 13'h0754
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_12_ERR_INTRO_Q0_1_12_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_12_ERR_INTRO_Q0_1_12_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_12_ERR_INTRO_Q0_1_12_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_12_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_12_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_12_BYTE_OFFSET 13'h0758
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_13_ERR_INTRO_Q0_1_13_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_13_ERR_INTRO_Q0_1_13_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_13_ERR_INTRO_Q0_1_13_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_13_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_13_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_13_BYTE_OFFSET 13'h075c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_14_ERR_INTRO_Q0_1_14_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_14_ERR_INTRO_Q0_1_14_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_14_ERR_INTRO_Q0_1_14_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_14_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_14_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_14_BYTE_OFFSET 13'h0760
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_15_ERR_INTRO_Q0_1_15_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_15_ERR_INTRO_Q0_1_15_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_15_ERR_INTRO_Q0_1_15_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_15_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_15_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_15_BYTE_OFFSET 13'h0764
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_16_ERR_INTRO_Q0_1_16_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_16_ERR_INTRO_Q0_1_16_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_16_ERR_INTRO_Q0_1_16_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_16_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_16_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_16_BYTE_OFFSET 13'h0768
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_17_ERR_INTRO_Q0_1_17_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_17_ERR_INTRO_Q0_1_17_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_17_ERR_INTRO_Q0_1_17_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_17_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_17_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_17_BYTE_OFFSET 13'h076c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_18_ERR_INTRO_Q0_1_18_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_18_ERR_INTRO_Q0_1_18_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_18_ERR_INTRO_Q0_1_18_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_18_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_18_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_18_BYTE_OFFSET 13'h0770
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_19_ERR_INTRO_Q0_1_19_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_19_ERR_INTRO_Q0_1_19_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_19_ERR_INTRO_Q0_1_19_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_19_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_19_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_19_BYTE_OFFSET 13'h0774
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_20_ERR_INTRO_Q0_1_20_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_20_ERR_INTRO_Q0_1_20_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_20_ERR_INTRO_Q0_1_20_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_20_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_20_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_20_BYTE_OFFSET 13'h0778
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_21_ERR_INTRO_Q0_1_21_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_21_ERR_INTRO_Q0_1_21_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_21_ERR_INTRO_Q0_1_21_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_21_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_21_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_21_BYTE_OFFSET 13'h077c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_22_ERR_INTRO_Q0_1_22_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_22_ERR_INTRO_Q0_1_22_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_22_ERR_INTRO_Q0_1_22_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_22_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_22_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_22_BYTE_OFFSET 13'h0780
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_23_ERR_INTRO_Q0_1_23_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_23_ERR_INTRO_Q0_1_23_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_23_ERR_INTRO_Q0_1_23_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_23_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_23_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_23_BYTE_OFFSET 13'h0784
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_24_ERR_INTRO_Q0_1_24_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_24_ERR_INTRO_Q0_1_24_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_24_ERR_INTRO_Q0_1_24_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_24_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_24_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_24_BYTE_OFFSET 13'h0788
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_25_ERR_INTRO_Q0_1_25_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_25_ERR_INTRO_Q0_1_25_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_25_ERR_INTRO_Q0_1_25_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_25_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_25_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_25_BYTE_OFFSET 13'h078c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_26_ERR_INTRO_Q0_1_26_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_26_ERR_INTRO_Q0_1_26_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_26_ERR_INTRO_Q0_1_26_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_26_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_26_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_26_BYTE_OFFSET 13'h0790
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_27_ERR_INTRO_Q0_1_27_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_27_ERR_INTRO_Q0_1_27_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_27_ERR_INTRO_Q0_1_27_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_27_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_27_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_27_BYTE_OFFSET 13'h0794
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_28_ERR_INTRO_Q0_1_28_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_28_ERR_INTRO_Q0_1_28_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_28_ERR_INTRO_Q0_1_28_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_28_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_28_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_28_BYTE_OFFSET 13'h0798
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_29_ERR_INTRO_Q0_1_29_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_29_ERR_INTRO_Q0_1_29_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_29_ERR_INTRO_Q0_1_29_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_29_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_29_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_29_BYTE_OFFSET 13'h079c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_30_ERR_INTRO_Q0_1_30_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_30_ERR_INTRO_Q0_1_30_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_30_ERR_INTRO_Q0_1_30_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_30_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_30_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_30_BYTE_OFFSET 13'h07a0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_31_ERR_INTRO_Q0_1_31_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_31_ERR_INTRO_Q0_1_31_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_31_ERR_INTRO_Q0_1_31_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_31_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_31_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_31_BYTE_OFFSET 13'h07a4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_32_ERR_INTRO_Q0_1_32_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_32_ERR_INTRO_Q0_1_32_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_32_ERR_INTRO_Q0_1_32_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_32_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_32_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_32_BYTE_OFFSET 13'h07a8
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_33_ERR_INTRO_Q0_1_33_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_33_ERR_INTRO_Q0_1_33_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_33_ERR_INTRO_Q0_1_33_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_33_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_33_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_33_BYTE_OFFSET 13'h07ac
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_34_ERR_INTRO_Q0_1_34_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_34_ERR_INTRO_Q0_1_34_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_34_ERR_INTRO_Q0_1_34_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_34_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_34_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_34_BYTE_OFFSET 13'h07b0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_35_ERR_INTRO_Q0_1_35_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_35_ERR_INTRO_Q0_1_35_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_35_ERR_INTRO_Q0_1_35_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_35_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_35_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_35_BYTE_OFFSET 13'h07b4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_36_ERR_INTRO_Q0_1_36_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_36_ERR_INTRO_Q0_1_36_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_36_ERR_INTRO_Q0_1_36_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_36_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_36_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_36_BYTE_OFFSET 13'h07b8
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_37_ERR_INTRO_Q0_1_37_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_37_ERR_INTRO_Q0_1_37_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_37_ERR_INTRO_Q0_1_37_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_37_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_37_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_37_BYTE_OFFSET 13'h07bc
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_38_ERR_INTRO_Q0_1_38_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_38_ERR_INTRO_Q0_1_38_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_38_ERR_INTRO_Q0_1_38_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_38_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_38_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_38_BYTE_OFFSET 13'h07c0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_39_ERR_INTRO_Q0_1_39_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_39_ERR_INTRO_Q0_1_39_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_39_ERR_INTRO_Q0_1_39_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_39_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_39_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_39_BYTE_OFFSET 13'h07c4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_40_ERR_INTRO_Q0_1_40_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_40_ERR_INTRO_Q0_1_40_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_40_ERR_INTRO_Q0_1_40_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_40_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_40_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_40_BYTE_OFFSET 13'h07c8
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_41_ERR_INTRO_Q0_1_41_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_41_ERR_INTRO_Q0_1_41_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_41_ERR_INTRO_Q0_1_41_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_41_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_41_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_41_BYTE_OFFSET 13'h07cc
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_42_ERR_INTRO_Q0_1_42_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_42_ERR_INTRO_Q0_1_42_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_42_ERR_INTRO_Q0_1_42_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_42_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_42_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_42_BYTE_OFFSET 13'h07d0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_43_ERR_INTRO_Q0_1_43_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_43_ERR_INTRO_Q0_1_43_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_43_ERR_INTRO_Q0_1_43_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_43_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_43_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_43_BYTE_OFFSET 13'h07d4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_44_ERR_INTRO_Q0_1_44_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_44_ERR_INTRO_Q0_1_44_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_44_ERR_INTRO_Q0_1_44_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_44_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_44_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_44_BYTE_OFFSET 13'h07d8
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_45_ERR_INTRO_Q0_1_45_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_45_ERR_INTRO_Q0_1_45_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_45_ERR_INTRO_Q0_1_45_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_45_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_45_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_45_BYTE_OFFSET 13'h07dc
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_46_ERR_INTRO_Q0_1_46_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_46_ERR_INTRO_Q0_1_46_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_46_ERR_INTRO_Q0_1_46_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_46_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_46_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_46_BYTE_OFFSET 13'h07e0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_47_ERR_INTRO_Q0_1_47_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_47_ERR_INTRO_Q0_1_47_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_47_ERR_INTRO_Q0_1_47_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_47_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_47_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_47_BYTE_OFFSET 13'h07e4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_48_ERR_INTRO_Q0_1_48_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_48_ERR_INTRO_Q0_1_48_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_48_ERR_INTRO_Q0_1_48_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_48_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_48_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_48_BYTE_OFFSET 13'h07e8
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_49_ERR_INTRO_Q0_1_49_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_49_ERR_INTRO_Q0_1_49_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_49_ERR_INTRO_Q0_1_49_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_49_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_49_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_49_BYTE_OFFSET 13'h07ec
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_50_ERR_INTRO_Q0_1_50_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_50_ERR_INTRO_Q0_1_50_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_50_ERR_INTRO_Q0_1_50_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_50_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_50_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_50_BYTE_OFFSET 13'h07f0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_51_ERR_INTRO_Q0_1_51_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_51_ERR_INTRO_Q0_1_51_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_51_ERR_INTRO_Q0_1_51_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_51_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_51_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_51_BYTE_OFFSET 13'h07f4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_52_ERR_INTRO_Q0_1_52_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_52_ERR_INTRO_Q0_1_52_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_52_ERR_INTRO_Q0_1_52_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_52_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_52_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_52_BYTE_OFFSET 13'h07f8
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_53_ERR_INTRO_Q0_1_53_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_53_ERR_INTRO_Q0_1_53_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_53_ERR_INTRO_Q0_1_53_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_53_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_53_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_53_BYTE_OFFSET 13'h07fc
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_54_ERR_INTRO_Q0_1_54_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_54_ERR_INTRO_Q0_1_54_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_54_ERR_INTRO_Q0_1_54_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_54_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_54_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_54_BYTE_OFFSET 13'h0800
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_55_ERR_INTRO_Q0_1_55_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_55_ERR_INTRO_Q0_1_55_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_55_ERR_INTRO_Q0_1_55_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_55_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_55_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_55_BYTE_OFFSET 13'h0804
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_56_ERR_INTRO_Q0_1_56_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_56_ERR_INTRO_Q0_1_56_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_56_ERR_INTRO_Q0_1_56_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_56_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_56_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_56_BYTE_OFFSET 13'h0808
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_57_ERR_INTRO_Q0_1_57_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_57_ERR_INTRO_Q0_1_57_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_57_ERR_INTRO_Q0_1_57_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_57_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_57_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_57_BYTE_OFFSET 13'h080c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_58_ERR_INTRO_Q0_1_58_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_58_ERR_INTRO_Q0_1_58_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_58_ERR_INTRO_Q0_1_58_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_58_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_58_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_58_BYTE_OFFSET 13'h0810
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_59_ERR_INTRO_Q0_1_59_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_59_ERR_INTRO_Q0_1_59_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_59_ERR_INTRO_Q0_1_59_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_59_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_59_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_59_BYTE_OFFSET 13'h0814
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_60_ERR_INTRO_Q0_1_60_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_60_ERR_INTRO_Q0_1_60_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_60_ERR_INTRO_Q0_1_60_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_60_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_60_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_60_BYTE_OFFSET 13'h0818
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_61_ERR_INTRO_Q0_1_61_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_61_ERR_INTRO_Q0_1_61_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_61_ERR_INTRO_Q0_1_61_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_61_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_61_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_61_BYTE_OFFSET 13'h081c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_62_ERR_INTRO_Q0_1_62_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_62_ERR_INTRO_Q0_1_62_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_62_ERR_INTRO_Q0_1_62_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_62_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_62_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_62_BYTE_OFFSET 13'h0820
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_63_ERR_INTRO_Q0_1_63_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_63_ERR_INTRO_Q0_1_63_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_63_ERR_INTRO_Q0_1_63_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_63_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_63_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_63_BYTE_OFFSET 13'h0824
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_64_ERR_INTRO_Q0_1_64_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_64_ERR_INTRO_Q0_1_64_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_64_ERR_INTRO_Q0_1_64_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_64_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_64_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_64_BYTE_OFFSET 13'h0828
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_65_ERR_INTRO_Q0_1_65_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_65_ERR_INTRO_Q0_1_65_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_65_ERR_INTRO_Q0_1_65_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_65_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_65_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_65_BYTE_OFFSET 13'h082c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_66_ERR_INTRO_Q0_1_66_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_66_ERR_INTRO_Q0_1_66_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_66_ERR_INTRO_Q0_1_66_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_66_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_66_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_66_BYTE_OFFSET 13'h0830
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_67_ERR_INTRO_Q0_1_67_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_67_ERR_INTRO_Q0_1_67_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_67_ERR_INTRO_Q0_1_67_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_67_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_67_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_67_BYTE_OFFSET 13'h0834
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_68_ERR_INTRO_Q0_1_68_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_68_ERR_INTRO_Q0_1_68_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_68_ERR_INTRO_Q0_1_68_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_68_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_68_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_68_BYTE_OFFSET 13'h0838
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_69_ERR_INTRO_Q0_1_69_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_69_ERR_INTRO_Q0_1_69_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_69_ERR_INTRO_Q0_1_69_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_69_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_69_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_69_BYTE_OFFSET 13'h083c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_70_ERR_INTRO_Q0_1_70_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_70_ERR_INTRO_Q0_1_70_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_70_ERR_INTRO_Q0_1_70_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_70_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_70_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_70_BYTE_OFFSET 13'h0840
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_71_ERR_INTRO_Q0_1_71_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_71_ERR_INTRO_Q0_1_71_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_71_ERR_INTRO_Q0_1_71_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_71_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_71_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_71_BYTE_OFFSET 13'h0844
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_72_ERR_INTRO_Q0_1_72_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_72_ERR_INTRO_Q0_1_72_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_72_ERR_INTRO_Q0_1_72_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_72_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_72_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_72_BYTE_OFFSET 13'h0848
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_73_ERR_INTRO_Q0_1_73_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_73_ERR_INTRO_Q0_1_73_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_73_ERR_INTRO_Q0_1_73_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_73_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_73_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_73_BYTE_OFFSET 13'h084c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_74_ERR_INTRO_Q0_1_74_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_74_ERR_INTRO_Q0_1_74_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_74_ERR_INTRO_Q0_1_74_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_74_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_74_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_74_BYTE_OFFSET 13'h0850
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_75_ERR_INTRO_Q0_1_75_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_75_ERR_INTRO_Q0_1_75_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_75_ERR_INTRO_Q0_1_75_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_75_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_75_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_75_BYTE_OFFSET 13'h0854
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_76_ERR_INTRO_Q0_1_76_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_76_ERR_INTRO_Q0_1_76_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_76_ERR_INTRO_Q0_1_76_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_76_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_76_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_76_BYTE_OFFSET 13'h0858
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_77_ERR_INTRO_Q0_1_77_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_77_ERR_INTRO_Q0_1_77_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_77_ERR_INTRO_Q0_1_77_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_77_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_77_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_77_BYTE_OFFSET 13'h085c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_78_ERR_INTRO_Q0_1_78_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_78_ERR_INTRO_Q0_1_78_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_78_ERR_INTRO_Q0_1_78_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_78_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_78_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_78_BYTE_OFFSET 13'h0860
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_79_ERR_INTRO_Q0_1_79_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_79_ERR_INTRO_Q0_1_79_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_79_ERR_INTRO_Q0_1_79_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_79_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_79_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_79_BYTE_OFFSET 13'h0864
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_80_ERR_INTRO_Q0_1_80_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_80_ERR_INTRO_Q0_1_80_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_80_ERR_INTRO_Q0_1_80_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_80_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_80_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_80_BYTE_OFFSET 13'h0868
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_81_ERR_INTRO_Q0_1_81_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_81_ERR_INTRO_Q0_1_81_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_81_ERR_INTRO_Q0_1_81_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_81_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_81_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_81_BYTE_OFFSET 13'h086c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_82_ERR_INTRO_Q0_1_82_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_82_ERR_INTRO_Q0_1_82_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_82_ERR_INTRO_Q0_1_82_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_82_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_82_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_82_BYTE_OFFSET 13'h0870
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_83_ERR_INTRO_Q0_1_83_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_83_ERR_INTRO_Q0_1_83_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_83_ERR_INTRO_Q0_1_83_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_83_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_83_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_83_BYTE_OFFSET 13'h0874
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_84_ERR_INTRO_Q0_1_84_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_84_ERR_INTRO_Q0_1_84_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_84_ERR_INTRO_Q0_1_84_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_84_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_84_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_84_BYTE_OFFSET 13'h0878
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_85_ERR_INTRO_Q0_1_85_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_85_ERR_INTRO_Q0_1_85_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_85_ERR_INTRO_Q0_1_85_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_85_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_85_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_85_BYTE_OFFSET 13'h087c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_86_ERR_INTRO_Q0_1_86_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_86_ERR_INTRO_Q0_1_86_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_86_ERR_INTRO_Q0_1_86_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_86_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_86_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_86_BYTE_OFFSET 13'h0880
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_87_ERR_INTRO_Q0_1_87_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_87_ERR_INTRO_Q0_1_87_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_87_ERR_INTRO_Q0_1_87_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_87_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_87_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_87_BYTE_OFFSET 13'h0884
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_88_ERR_INTRO_Q0_1_88_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_88_ERR_INTRO_Q0_1_88_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_88_ERR_INTRO_Q0_1_88_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_88_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_88_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_88_BYTE_OFFSET 13'h0888
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_89_ERR_INTRO_Q0_1_89_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_89_ERR_INTRO_Q0_1_89_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_89_ERR_INTRO_Q0_1_89_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_89_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_89_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_89_BYTE_OFFSET 13'h088c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_90_ERR_INTRO_Q0_1_90_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_90_ERR_INTRO_Q0_1_90_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_90_ERR_INTRO_Q0_1_90_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_90_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_90_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_90_BYTE_OFFSET 13'h0890
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_91_ERR_INTRO_Q0_1_91_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_91_ERR_INTRO_Q0_1_91_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_91_ERR_INTRO_Q0_1_91_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_91_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_91_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_91_BYTE_OFFSET 13'h0894
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_92_ERR_INTRO_Q0_1_92_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_92_ERR_INTRO_Q0_1_92_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_92_ERR_INTRO_Q0_1_92_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_92_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_92_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_92_BYTE_OFFSET 13'h0898
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_93_ERR_INTRO_Q0_1_93_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_93_ERR_INTRO_Q0_1_93_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_93_ERR_INTRO_Q0_1_93_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_93_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_93_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_93_BYTE_OFFSET 13'h089c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_94_ERR_INTRO_Q0_1_94_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_94_ERR_INTRO_Q0_1_94_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_94_ERR_INTRO_Q0_1_94_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_94_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_94_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_94_BYTE_OFFSET 13'h08a0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_95_ERR_INTRO_Q0_1_95_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_95_ERR_INTRO_Q0_1_95_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_95_ERR_INTRO_Q0_1_95_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_95_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_95_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_95_BYTE_OFFSET 13'h08a4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_96_ERR_INTRO_Q0_1_96_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_96_ERR_INTRO_Q0_1_96_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_96_ERR_INTRO_Q0_1_96_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_96_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_96_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_96_BYTE_OFFSET 13'h08a8
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_97_ERR_INTRO_Q0_1_97_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_97_ERR_INTRO_Q0_1_97_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_97_ERR_INTRO_Q0_1_97_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_97_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_97_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_97_BYTE_OFFSET 13'h08ac
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_98_ERR_INTRO_Q0_1_98_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_98_ERR_INTRO_Q0_1_98_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_98_ERR_INTRO_Q0_1_98_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_98_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_98_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_98_BYTE_OFFSET 13'h08b0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_99_ERR_INTRO_Q0_1_99_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_99_ERR_INTRO_Q0_1_99_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_99_ERR_INTRO_Q0_1_99_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_99_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_99_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_99_BYTE_OFFSET 13'h08b4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_100_ERR_INTRO_Q0_1_100_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_100_ERR_INTRO_Q0_1_100_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_100_ERR_INTRO_Q0_1_100_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_100_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_100_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_100_BYTE_OFFSET 13'h08b8
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_101_ERR_INTRO_Q0_1_101_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_101_ERR_INTRO_Q0_1_101_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_101_ERR_INTRO_Q0_1_101_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_101_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_101_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_101_BYTE_OFFSET 13'h08bc
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_102_ERR_INTRO_Q0_1_102_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_102_ERR_INTRO_Q0_1_102_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_102_ERR_INTRO_Q0_1_102_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_102_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_102_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_102_BYTE_OFFSET 13'h08c0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_103_ERR_INTRO_Q0_1_103_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_103_ERR_INTRO_Q0_1_103_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_103_ERR_INTRO_Q0_1_103_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_103_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_103_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_103_BYTE_OFFSET 13'h08c4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_104_ERR_INTRO_Q0_1_104_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_104_ERR_INTRO_Q0_1_104_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_104_ERR_INTRO_Q0_1_104_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_104_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_104_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_104_BYTE_OFFSET 13'h08c8
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_105_ERR_INTRO_Q0_1_105_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_105_ERR_INTRO_Q0_1_105_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_105_ERR_INTRO_Q0_1_105_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_105_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_105_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_105_BYTE_OFFSET 13'h08cc
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_106_ERR_INTRO_Q0_1_106_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_106_ERR_INTRO_Q0_1_106_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_106_ERR_INTRO_Q0_1_106_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_106_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_106_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_106_BYTE_OFFSET 13'h08d0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_107_ERR_INTRO_Q0_1_107_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_107_ERR_INTRO_Q0_1_107_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_107_ERR_INTRO_Q0_1_107_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_107_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_107_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_107_BYTE_OFFSET 13'h08d4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_108_ERR_INTRO_Q0_1_108_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_108_ERR_INTRO_Q0_1_108_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_108_ERR_INTRO_Q0_1_108_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_108_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_108_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_108_BYTE_OFFSET 13'h08d8
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_109_ERR_INTRO_Q0_1_109_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_109_ERR_INTRO_Q0_1_109_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_109_ERR_INTRO_Q0_1_109_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_109_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_109_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_109_BYTE_OFFSET 13'h08dc
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_110_ERR_INTRO_Q0_1_110_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_110_ERR_INTRO_Q0_1_110_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_110_ERR_INTRO_Q0_1_110_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_110_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_110_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_110_BYTE_OFFSET 13'h08e0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_111_ERR_INTRO_Q0_1_111_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_111_ERR_INTRO_Q0_1_111_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_111_ERR_INTRO_Q0_1_111_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_111_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_111_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_111_BYTE_OFFSET 13'h08e4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_112_ERR_INTRO_Q0_1_112_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_112_ERR_INTRO_Q0_1_112_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_112_ERR_INTRO_Q0_1_112_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_112_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_112_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_112_BYTE_OFFSET 13'h08e8
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_113_ERR_INTRO_Q0_1_113_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_113_ERR_INTRO_Q0_1_113_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_113_ERR_INTRO_Q0_1_113_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_113_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_113_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_113_BYTE_OFFSET 13'h08ec
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_114_ERR_INTRO_Q0_1_114_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_114_ERR_INTRO_Q0_1_114_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_114_ERR_INTRO_Q0_1_114_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_114_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_114_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_114_BYTE_OFFSET 13'h08f0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_115_ERR_INTRO_Q0_1_115_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_115_ERR_INTRO_Q0_1_115_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_115_ERR_INTRO_Q0_1_115_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_115_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_115_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_115_BYTE_OFFSET 13'h08f4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_116_ERR_INTRO_Q0_1_116_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_116_ERR_INTRO_Q0_1_116_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_116_ERR_INTRO_Q0_1_116_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_116_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_116_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_116_BYTE_OFFSET 13'h08f8
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_117_ERR_INTRO_Q0_1_117_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_117_ERR_INTRO_Q0_1_117_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_117_ERR_INTRO_Q0_1_117_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_117_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_117_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_117_BYTE_OFFSET 13'h08fc
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_118_ERR_INTRO_Q0_1_118_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_118_ERR_INTRO_Q0_1_118_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_118_ERR_INTRO_Q0_1_118_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_118_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_118_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_118_BYTE_OFFSET 13'h0900
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_119_ERR_INTRO_Q0_1_119_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_119_ERR_INTRO_Q0_1_119_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_119_ERR_INTRO_Q0_1_119_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_119_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_119_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_119_BYTE_OFFSET 13'h0904
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_120_ERR_INTRO_Q0_1_120_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_120_ERR_INTRO_Q0_1_120_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_120_ERR_INTRO_Q0_1_120_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_120_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_120_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_120_BYTE_OFFSET 13'h0908
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_121_ERR_INTRO_Q0_1_121_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_121_ERR_INTRO_Q0_1_121_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_121_ERR_INTRO_Q0_1_121_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_121_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_121_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_121_BYTE_OFFSET 13'h090c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_122_ERR_INTRO_Q0_1_122_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_122_ERR_INTRO_Q0_1_122_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_122_ERR_INTRO_Q0_1_122_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_122_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_122_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_122_BYTE_OFFSET 13'h0910
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_123_ERR_INTRO_Q0_1_123_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_123_ERR_INTRO_Q0_1_123_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_123_ERR_INTRO_Q0_1_123_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_123_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_123_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_123_BYTE_OFFSET 13'h0914
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_124_ERR_INTRO_Q0_1_124_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_124_ERR_INTRO_Q0_1_124_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_124_ERR_INTRO_Q0_1_124_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_124_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_124_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_124_BYTE_OFFSET 13'h0918
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_125_ERR_INTRO_Q0_1_125_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_125_ERR_INTRO_Q0_1_125_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_125_ERR_INTRO_Q0_1_125_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_125_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_125_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_125_BYTE_OFFSET 13'h091c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_126_ERR_INTRO_Q0_1_126_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_126_ERR_INTRO_Q0_1_126_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_126_ERR_INTRO_Q0_1_126_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_126_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_126_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_126_BYTE_OFFSET 13'h0920
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_127_ERR_INTRO_Q0_1_127_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_127_ERR_INTRO_Q0_1_127_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_127_ERR_INTRO_Q0_1_127_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_127_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_127_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_127_BYTE_OFFSET 13'h0924
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_128_ERR_INTRO_Q0_1_128_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_128_ERR_INTRO_Q0_1_128_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_128_ERR_INTRO_Q0_1_128_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_128_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_128_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_128_BYTE_OFFSET 13'h0928
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_129_ERR_INTRO_Q0_1_129_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_129_ERR_INTRO_Q0_1_129_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_129_ERR_INTRO_Q0_1_129_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_129_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_129_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_129_BYTE_OFFSET 13'h092c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_130_ERR_INTRO_Q0_1_130_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_130_ERR_INTRO_Q0_1_130_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_130_ERR_INTRO_Q0_1_130_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_130_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_130_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_130_BYTE_OFFSET 13'h0930
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_131_ERR_INTRO_Q0_1_131_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_131_ERR_INTRO_Q0_1_131_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_131_ERR_INTRO_Q0_1_131_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_131_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_131_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_131_BYTE_OFFSET 13'h0934
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_132_ERR_INTRO_Q0_1_132_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_132_ERR_INTRO_Q0_1_132_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_132_ERR_INTRO_Q0_1_132_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_132_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_132_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_132_BYTE_OFFSET 13'h0938
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_133_ERR_INTRO_Q0_1_133_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_133_ERR_INTRO_Q0_1_133_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_133_ERR_INTRO_Q0_1_133_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_133_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_133_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_133_BYTE_OFFSET 13'h093c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_134_ERR_INTRO_Q0_1_134_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_134_ERR_INTRO_Q0_1_134_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_134_ERR_INTRO_Q0_1_134_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_134_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_134_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_134_BYTE_OFFSET 13'h0940
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_135_ERR_INTRO_Q0_1_135_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_135_ERR_INTRO_Q0_1_135_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_135_ERR_INTRO_Q0_1_135_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_135_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_135_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_135_BYTE_OFFSET 13'h0944
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_136_ERR_INTRO_Q0_1_136_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_136_ERR_INTRO_Q0_1_136_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_136_ERR_INTRO_Q0_1_136_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_136_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_136_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_136_BYTE_OFFSET 13'h0948
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_137_ERR_INTRO_Q0_1_137_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_137_ERR_INTRO_Q0_1_137_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_137_ERR_INTRO_Q0_1_137_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_137_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_137_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_137_BYTE_OFFSET 13'h094c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_138_ERR_INTRO_Q0_1_138_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_138_ERR_INTRO_Q0_1_138_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_138_ERR_INTRO_Q0_1_138_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_138_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_138_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_138_BYTE_OFFSET 13'h0950
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_139_ERR_INTRO_Q0_1_139_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_139_ERR_INTRO_Q0_1_139_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_139_ERR_INTRO_Q0_1_139_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_139_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_139_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_139_BYTE_OFFSET 13'h0954
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_140_ERR_INTRO_Q0_1_140_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_140_ERR_INTRO_Q0_1_140_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_140_ERR_INTRO_Q0_1_140_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_140_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_140_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_140_BYTE_OFFSET 13'h0958
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_141_ERR_INTRO_Q0_1_141_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_141_ERR_INTRO_Q0_1_141_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_141_ERR_INTRO_Q0_1_141_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_141_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_141_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_141_BYTE_OFFSET 13'h095c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_142_ERR_INTRO_Q0_1_142_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_142_ERR_INTRO_Q0_1_142_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_142_ERR_INTRO_Q0_1_142_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_142_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_142_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_142_BYTE_OFFSET 13'h0960
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_143_ERR_INTRO_Q0_1_143_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_143_ERR_INTRO_Q0_1_143_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_143_ERR_INTRO_Q0_1_143_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_143_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_143_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_143_BYTE_OFFSET 13'h0964
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_144_ERR_INTRO_Q0_1_144_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_144_ERR_INTRO_Q0_1_144_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_144_ERR_INTRO_Q0_1_144_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_144_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_144_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_144_BYTE_OFFSET 13'h0968
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_145_ERR_INTRO_Q0_1_145_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_145_ERR_INTRO_Q0_1_145_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_145_ERR_INTRO_Q0_1_145_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_145_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_145_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_145_BYTE_OFFSET 13'h096c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_146_ERR_INTRO_Q0_1_146_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_146_ERR_INTRO_Q0_1_146_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_146_ERR_INTRO_Q0_1_146_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_146_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_146_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_146_BYTE_OFFSET 13'h0970
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_147_ERR_INTRO_Q0_1_147_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_147_ERR_INTRO_Q0_1_147_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_147_ERR_INTRO_Q0_1_147_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_147_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_147_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_147_BYTE_OFFSET 13'h0974
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_148_ERR_INTRO_Q0_1_148_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_148_ERR_INTRO_Q0_1_148_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_148_ERR_INTRO_Q0_1_148_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_148_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_148_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_148_BYTE_OFFSET 13'h0978
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_149_ERR_INTRO_Q0_1_149_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_149_ERR_INTRO_Q0_1_149_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_149_ERR_INTRO_Q0_1_149_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_149_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_149_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_149_BYTE_OFFSET 13'h097c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_150_ERR_INTRO_Q0_1_150_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_150_ERR_INTRO_Q0_1_150_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_150_ERR_INTRO_Q0_1_150_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_150_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_150_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_150_BYTE_OFFSET 13'h0980
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_151_ERR_INTRO_Q0_1_151_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_151_ERR_INTRO_Q0_1_151_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_151_ERR_INTRO_Q0_1_151_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_151_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_151_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_151_BYTE_OFFSET 13'h0984
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_152_ERR_INTRO_Q0_1_152_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_152_ERR_INTRO_Q0_1_152_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_152_ERR_INTRO_Q0_1_152_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_152_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_152_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_152_BYTE_OFFSET 13'h0988
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_153_ERR_INTRO_Q0_1_153_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_153_ERR_INTRO_Q0_1_153_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_153_ERR_INTRO_Q0_1_153_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_153_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_153_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_153_BYTE_OFFSET 13'h098c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_154_ERR_INTRO_Q0_1_154_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_154_ERR_INTRO_Q0_1_154_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_154_ERR_INTRO_Q0_1_154_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_154_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_154_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_154_BYTE_OFFSET 13'h0990
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_155_ERR_INTRO_Q0_1_155_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_155_ERR_INTRO_Q0_1_155_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_155_ERR_INTRO_Q0_1_155_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_155_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_155_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_155_BYTE_OFFSET 13'h0994
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_156_ERR_INTRO_Q0_1_156_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_156_ERR_INTRO_Q0_1_156_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_156_ERR_INTRO_Q0_1_156_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_156_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_156_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_156_BYTE_OFFSET 13'h0998
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_157_ERR_INTRO_Q0_1_157_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_157_ERR_INTRO_Q0_1_157_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_157_ERR_INTRO_Q0_1_157_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_157_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_157_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_157_BYTE_OFFSET 13'h099c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_158_ERR_INTRO_Q0_1_158_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_158_ERR_INTRO_Q0_1_158_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_158_ERR_INTRO_Q0_1_158_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_158_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_158_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_158_BYTE_OFFSET 13'h09a0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_159_ERR_INTRO_Q0_1_159_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_159_ERR_INTRO_Q0_1_159_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_159_ERR_INTRO_Q0_1_159_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_159_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_159_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_159_BYTE_OFFSET 13'h09a4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_160_ERR_INTRO_Q0_1_160_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_160_ERR_INTRO_Q0_1_160_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_160_ERR_INTRO_Q0_1_160_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_160_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_160_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_160_BYTE_OFFSET 13'h09a8
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_161_ERR_INTRO_Q0_1_161_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_161_ERR_INTRO_Q0_1_161_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_161_ERR_INTRO_Q0_1_161_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_161_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_161_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_161_BYTE_OFFSET 13'h09ac
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_162_ERR_INTRO_Q0_1_162_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_162_ERR_INTRO_Q0_1_162_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_162_ERR_INTRO_Q0_1_162_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_162_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_162_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_162_BYTE_OFFSET 13'h09b0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_163_ERR_INTRO_Q0_1_163_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_163_ERR_INTRO_Q0_1_163_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_163_ERR_INTRO_Q0_1_163_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_163_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_163_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_163_BYTE_OFFSET 13'h09b4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_164_ERR_INTRO_Q0_1_164_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_164_ERR_INTRO_Q0_1_164_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_164_ERR_INTRO_Q0_1_164_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_164_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_164_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_164_BYTE_OFFSET 13'h09b8
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_165_ERR_INTRO_Q0_1_165_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_165_ERR_INTRO_Q0_1_165_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_165_ERR_INTRO_Q0_1_165_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_165_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_165_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_165_BYTE_OFFSET 13'h09bc
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_166_ERR_INTRO_Q0_1_166_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_166_ERR_INTRO_Q0_1_166_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_166_ERR_INTRO_Q0_1_166_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_166_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_166_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_166_BYTE_OFFSET 13'h09c0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_167_ERR_INTRO_Q0_1_167_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_167_ERR_INTRO_Q0_1_167_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_167_ERR_INTRO_Q0_1_167_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_167_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_167_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_167_BYTE_OFFSET 13'h09c4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_168_ERR_INTRO_Q0_1_168_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_168_ERR_INTRO_Q0_1_168_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_168_ERR_INTRO_Q0_1_168_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_168_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_168_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_168_BYTE_OFFSET 13'h09c8
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_169_ERR_INTRO_Q0_1_169_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_169_ERR_INTRO_Q0_1_169_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_169_ERR_INTRO_Q0_1_169_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_169_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_169_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_169_BYTE_OFFSET 13'h09cc
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_170_ERR_INTRO_Q0_1_170_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_170_ERR_INTRO_Q0_1_170_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_170_ERR_INTRO_Q0_1_170_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_170_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_170_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_170_BYTE_OFFSET 13'h09d0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_171_ERR_INTRO_Q0_1_171_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_171_ERR_INTRO_Q0_1_171_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_171_ERR_INTRO_Q0_1_171_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_171_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_171_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_171_BYTE_OFFSET 13'h09d4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_172_ERR_INTRO_Q0_1_172_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_172_ERR_INTRO_Q0_1_172_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_172_ERR_INTRO_Q0_1_172_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_172_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_172_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_172_BYTE_OFFSET 13'h09d8
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_173_ERR_INTRO_Q0_1_173_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_173_ERR_INTRO_Q0_1_173_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_173_ERR_INTRO_Q0_1_173_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_173_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_173_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_173_BYTE_OFFSET 13'h09dc
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_174_ERR_INTRO_Q0_1_174_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_174_ERR_INTRO_Q0_1_174_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_174_ERR_INTRO_Q0_1_174_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_174_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_174_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_174_BYTE_OFFSET 13'h09e0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_175_ERR_INTRO_Q0_1_175_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_175_ERR_INTRO_Q0_1_175_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_175_ERR_INTRO_Q0_1_175_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_175_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_175_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_175_BYTE_OFFSET 13'h09e4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_176_ERR_INTRO_Q0_1_176_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_176_ERR_INTRO_Q0_1_176_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_176_ERR_INTRO_Q0_1_176_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_176_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_176_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_176_BYTE_OFFSET 13'h09e8
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_177_ERR_INTRO_Q0_1_177_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_177_ERR_INTRO_Q0_1_177_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_177_ERR_INTRO_Q0_1_177_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_177_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_177_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_177_BYTE_OFFSET 13'h09ec
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_178_ERR_INTRO_Q0_1_178_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_178_ERR_INTRO_Q0_1_178_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_178_ERR_INTRO_Q0_1_178_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_178_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_178_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_178_BYTE_OFFSET 13'h09f0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_179_ERR_INTRO_Q0_1_179_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_179_ERR_INTRO_Q0_1_179_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_179_ERR_INTRO_Q0_1_179_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_179_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_179_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_179_BYTE_OFFSET 13'h09f4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_180_ERR_INTRO_Q0_1_180_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_180_ERR_INTRO_Q0_1_180_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_180_ERR_INTRO_Q0_1_180_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_180_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_180_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_180_BYTE_OFFSET 13'h09f8
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_181_ERR_INTRO_Q0_1_181_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_181_ERR_INTRO_Q0_1_181_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_181_ERR_INTRO_Q0_1_181_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_181_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_181_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_181_BYTE_OFFSET 13'h09fc
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_182_ERR_INTRO_Q0_1_182_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_182_ERR_INTRO_Q0_1_182_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_182_ERR_INTRO_Q0_1_182_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_182_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_182_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_182_BYTE_OFFSET 13'h0a00
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_183_ERR_INTRO_Q0_1_183_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_183_ERR_INTRO_Q0_1_183_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_183_ERR_INTRO_Q0_1_183_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_183_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_183_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_183_BYTE_OFFSET 13'h0a04
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_184_ERR_INTRO_Q0_1_184_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_184_ERR_INTRO_Q0_1_184_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_184_ERR_INTRO_Q0_1_184_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_184_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_184_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_184_BYTE_OFFSET 13'h0a08
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_185_ERR_INTRO_Q0_1_185_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_185_ERR_INTRO_Q0_1_185_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_185_ERR_INTRO_Q0_1_185_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_185_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_185_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_185_BYTE_OFFSET 13'h0a0c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_186_ERR_INTRO_Q0_1_186_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_186_ERR_INTRO_Q0_1_186_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_186_ERR_INTRO_Q0_1_186_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_186_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_186_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_186_BYTE_OFFSET 13'h0a10
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_187_ERR_INTRO_Q0_1_187_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_187_ERR_INTRO_Q0_1_187_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_187_ERR_INTRO_Q0_1_187_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_187_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_187_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_187_BYTE_OFFSET 13'h0a14
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_188_ERR_INTRO_Q0_1_188_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_188_ERR_INTRO_Q0_1_188_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_188_ERR_INTRO_Q0_1_188_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_188_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_188_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_188_BYTE_OFFSET 13'h0a18
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_189_ERR_INTRO_Q0_1_189_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_189_ERR_INTRO_Q0_1_189_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_189_ERR_INTRO_Q0_1_189_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_189_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_189_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_189_BYTE_OFFSET 13'h0a1c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_190_ERR_INTRO_Q0_1_190_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_190_ERR_INTRO_Q0_1_190_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_190_ERR_INTRO_Q0_1_190_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_190_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_190_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_190_BYTE_OFFSET 13'h0a20
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_191_ERR_INTRO_Q0_1_191_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_191_ERR_INTRO_Q0_1_191_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_191_ERR_INTRO_Q0_1_191_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_191_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_191_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_191_BYTE_OFFSET 13'h0a24
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_192_ERR_INTRO_Q0_1_192_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_192_ERR_INTRO_Q0_1_192_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_192_ERR_INTRO_Q0_1_192_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_192_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_192_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_192_BYTE_OFFSET 13'h0a28
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_193_ERR_INTRO_Q0_1_193_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_193_ERR_INTRO_Q0_1_193_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_193_ERR_INTRO_Q0_1_193_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_193_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_193_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_193_BYTE_OFFSET 13'h0a2c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_194_ERR_INTRO_Q0_1_194_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_194_ERR_INTRO_Q0_1_194_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_194_ERR_INTRO_Q0_1_194_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_194_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_194_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_194_BYTE_OFFSET 13'h0a30
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_195_ERR_INTRO_Q0_1_195_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_195_ERR_INTRO_Q0_1_195_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_195_ERR_INTRO_Q0_1_195_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_195_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_195_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_195_BYTE_OFFSET 13'h0a34
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_196_ERR_INTRO_Q0_1_196_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_196_ERR_INTRO_Q0_1_196_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_196_ERR_INTRO_Q0_1_196_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_196_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_196_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_196_BYTE_OFFSET 13'h0a38
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_197_ERR_INTRO_Q0_1_197_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_197_ERR_INTRO_Q0_1_197_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_197_ERR_INTRO_Q0_1_197_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_197_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_197_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_197_BYTE_OFFSET 13'h0a3c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_198_ERR_INTRO_Q0_1_198_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_198_ERR_INTRO_Q0_1_198_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_198_ERR_INTRO_Q0_1_198_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_198_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_198_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_198_BYTE_OFFSET 13'h0a40
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_199_ERR_INTRO_Q0_1_199_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_199_ERR_INTRO_Q0_1_199_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_199_ERR_INTRO_Q0_1_199_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_199_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_199_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_199_BYTE_OFFSET 13'h0a44
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_200_ERR_INTRO_Q0_1_200_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_200_ERR_INTRO_Q0_1_200_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_200_ERR_INTRO_Q0_1_200_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_200_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_200_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_200_BYTE_OFFSET 13'h0a48
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_201_ERR_INTRO_Q0_1_201_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_201_ERR_INTRO_Q0_1_201_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_201_ERR_INTRO_Q0_1_201_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_201_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_201_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_201_BYTE_OFFSET 13'h0a4c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_202_ERR_INTRO_Q0_1_202_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_202_ERR_INTRO_Q0_1_202_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_202_ERR_INTRO_Q0_1_202_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_202_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_202_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_202_BYTE_OFFSET 13'h0a50
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_203_ERR_INTRO_Q0_1_203_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_203_ERR_INTRO_Q0_1_203_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_203_ERR_INTRO_Q0_1_203_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_203_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_203_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_203_BYTE_OFFSET 13'h0a54
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_204_ERR_INTRO_Q0_1_204_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_204_ERR_INTRO_Q0_1_204_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_204_ERR_INTRO_Q0_1_204_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_204_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_204_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_204_BYTE_OFFSET 13'h0a58
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_205_ERR_INTRO_Q0_1_205_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_205_ERR_INTRO_Q0_1_205_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_205_ERR_INTRO_Q0_1_205_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_205_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_205_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_205_BYTE_OFFSET 13'h0a5c
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_206_ERR_INTRO_Q0_1_206_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_206_ERR_INTRO_Q0_1_206_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_206_ERR_INTRO_Q0_1_206_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_206_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_206_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_206_BYTE_OFFSET 13'h0a60
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_207_ERR_INTRO_Q0_1_207_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_207_ERR_INTRO_Q0_1_207_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_207_ERR_INTRO_Q0_1_207_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_207_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_207_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_Q0_1_INTRO_207_BYTE_OFFSET 13'h0a64
`define LDPC_CSR_LDPC_DEC_ERR_INTRODUCED_ERR_INTRO_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_INTRODUCED_ERR_INTRO_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_INTRODUCED_ERR_INTRO_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_INTRODUCED_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_INTRODUCED_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_INTRODUCED_BYTE_OFFSET 13'h0a68
`define LDPC_CSR_LDPC_DEC_ERR_INTRO_DECODER_ERR_INTRO_DECODER_BIT_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_ERR_INTRO_DECODER_ERR_INTRO_DECODER_BIT_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_ERR_INTRO_DECODER_ERR_INTRO_DECODER_BIT_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_ERR_INTRO_DECODER_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_ERR_INTRO_DECODER_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_ERR_INTRO_DECODER_BYTE_OFFSET 13'h0a6c
`define LDPC_CSR_LDPC_DEC_PROBABILITY_PERC_PROBABILITY_BIT_WIDTH 32
`define LDPC_CSR_LDPC_DEC_PROBABILITY_PERC_PROBABILITY_BIT_MASK 32'hffffffff
`define LDPC_CSR_LDPC_DEC_PROBABILITY_PERC_PROBABILITY_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_PROBABILITY_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_PROBABILITY_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_PROBABILITY_BYTE_OFFSET 13'h0a70
`define LDPC_CSR_LDPC_DEC_HAMDIST_LOOP_MAX_HAMDIST_LOOP_MAX_BIT_WIDTH 32
`define LDPC_CSR_LDPC_DEC_HAMDIST_LOOP_MAX_HAMDIST_LOOP_MAX_BIT_MASK 32'hffffffff
`define LDPC_CSR_LDPC_DEC_HAMDIST_LOOP_MAX_HAMDIST_LOOP_MAX_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_HAMDIST_LOOP_MAX_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_HAMDIST_LOOP_MAX_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_HAMDIST_LOOP_MAX_BYTE_OFFSET 13'h0a74
`define LDPC_CSR_LDPC_DEC_HAMDIST_LOOP_PERCENTAGE_HAMDIST_LOOP_PERCENTAGE_BIT_WIDTH 32
`define LDPC_CSR_LDPC_DEC_HAMDIST_LOOP_PERCENTAGE_HAMDIST_LOOP_PERCENTAGE_BIT_MASK 32'hffffffff
`define LDPC_CSR_LDPC_DEC_HAMDIST_LOOP_PERCENTAGE_HAMDIST_LOOP_PERCENTAGE_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_HAMDIST_LOOP_PERCENTAGE_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_HAMDIST_LOOP_PERCENTAGE_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_HAMDIST_LOOP_PERCENTAGE_BYTE_OFFSET 13'h0a78
`define LDPC_CSR_LDPC_DEC_HAMDIST_IIR1_HAMDIST_IIR1_BIT_WIDTH 32
`define LDPC_CSR_LDPC_DEC_HAMDIST_IIR1_HAMDIST_IIR1_BIT_MASK 32'hffffffff
`define LDPC_CSR_LDPC_DEC_HAMDIST_IIR1_HAMDIST_IIR1_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_HAMDIST_IIR1_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_HAMDIST_IIR1_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_HAMDIST_IIR1_BYTE_OFFSET 13'h0a7c
`define LDPC_CSR_LDPC_DEC_HAMDIST_IIR2_NOT_USED_HAMDIST_IIR2_BIT_WIDTH 32
`define LDPC_CSR_LDPC_DEC_HAMDIST_IIR2_NOT_USED_HAMDIST_IIR2_BIT_MASK 32'hffffffff
`define LDPC_CSR_LDPC_DEC_HAMDIST_IIR2_NOT_USED_HAMDIST_IIR2_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_HAMDIST_IIR2_NOT_USED_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_HAMDIST_IIR2_NOT_USED_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_HAMDIST_IIR2_NOT_USED_BYTE_OFFSET 13'h0a80
`define LDPC_CSR_LDPC_DEC_HAMDIST_IIR3_NOT_USED_HAMDIST_IIR3_BIT_WIDTH 32
`define LDPC_CSR_LDPC_DEC_HAMDIST_IIR3_NOT_USED_HAMDIST_IIR3_BIT_MASK 32'hffffffff
`define LDPC_CSR_LDPC_DEC_HAMDIST_IIR3_NOT_USED_HAMDIST_IIR3_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_HAMDIST_IIR3_NOT_USED_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_HAMDIST_IIR3_NOT_USED_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_HAMDIST_IIR3_NOT_USED_BYTE_OFFSET 13'h0a84
`define LDPC_CSR_LDPC_DEC_SYN_VALID_CWORD_DEC_FINAL_SYN_VALID_CWORD_DEC_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_SYN_VALID_CWORD_DEC_FINAL_SYN_VALID_CWORD_DEC_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_SYN_VALID_CWORD_DEC_FINAL_SYN_VALID_CWORD_DEC_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_SYN_VALID_CWORD_DEC_FINAL_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_SYN_VALID_CWORD_DEC_FINAL_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_SYN_VALID_CWORD_DEC_FINAL_BYTE_OFFSET 13'h0a88
`define LDPC_CSR_LDPC_DEC_START_DEC_START_DEC_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_START_DEC_START_DEC_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_START_DEC_START_DEC_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_START_DEC_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_START_DEC_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_START_DEC_BYTE_OFFSET 13'h0a8c
`define LDPC_CSR_LDPC_DEC_CONVERGED_LOOPS_ENDED_CONVERGED_LOOPS_ENDED_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CONVERGED_LOOPS_ENDED_CONVERGED_LOOPS_ENDED_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CONVERGED_LOOPS_ENDED_CONVERGED_LOOPS_ENDED_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CONVERGED_LOOPS_ENDED_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CONVERGED_LOOPS_ENDED_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CONVERGED_LOOPS_ENDED_BYTE_OFFSET 13'h0a90
`define LDPC_CSR_LDPC_DEC_CONVERGED_PASS_FAIL_CONVERGED_PASS_FAIL_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CONVERGED_PASS_FAIL_CONVERGED_PASS_FAIL_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CONVERGED_PASS_FAIL_CONVERGED_PASS_FAIL_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CONVERGED_PASS_FAIL_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CONVERGED_PASS_FAIL_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CONVERGED_PASS_FAIL_BYTE_OFFSET 13'h0a94
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_0_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_0_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_0_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_0_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_0_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_0_BYTE_OFFSET 13'h0a98
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_1_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_1_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_1_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_1_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_1_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_1_BYTE_OFFSET 13'h0a9c
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_2_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_2_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_2_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_2_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_2_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_2_BYTE_OFFSET 13'h0aa0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_3_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_3_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_3_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_3_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_3_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_3_BYTE_OFFSET 13'h0aa4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_4_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_4_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_4_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_4_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_4_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_4_BYTE_OFFSET 13'h0aa8
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_5_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_5_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_5_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_5_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_5_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_5_BYTE_OFFSET 13'h0aac
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_6_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_6_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_6_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_6_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_6_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_6_BYTE_OFFSET 13'h0ab0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_7_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_7_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_7_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_7_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_7_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_7_BYTE_OFFSET 13'h0ab4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_8_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_8_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_8_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_8_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_8_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_8_BYTE_OFFSET 13'h0ab8
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_9_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_9_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_9_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_9_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_9_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_9_BYTE_OFFSET 13'h0abc
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_10_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_10_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_10_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_10_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_10_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_10_BYTE_OFFSET 13'h0ac0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_11_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_11_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_11_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_11_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_11_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_11_BYTE_OFFSET 13'h0ac4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_12_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_12_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_12_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_12_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_12_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_12_BYTE_OFFSET 13'h0ac8
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_13_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_13_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_13_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_13_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_13_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_13_BYTE_OFFSET 13'h0acc
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_14_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_14_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_14_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_14_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_14_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_14_BYTE_OFFSET 13'h0ad0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_15_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_15_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_15_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_15_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_15_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_15_BYTE_OFFSET 13'h0ad4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_16_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_16_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_16_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_16_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_16_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_16_BYTE_OFFSET 13'h0ad8
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_17_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_17_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_17_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_17_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_17_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_17_BYTE_OFFSET 13'h0adc
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_18_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_18_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_18_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_18_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_18_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_18_BYTE_OFFSET 13'h0ae0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_19_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_19_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_19_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_19_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_19_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_19_BYTE_OFFSET 13'h0ae4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_20_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_20_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_20_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_20_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_20_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_20_BYTE_OFFSET 13'h0ae8
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_21_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_21_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_21_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_21_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_21_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_21_BYTE_OFFSET 13'h0aec
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_22_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_22_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_22_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_22_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_22_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_22_BYTE_OFFSET 13'h0af0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_23_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_23_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_23_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_23_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_23_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_23_BYTE_OFFSET 13'h0af4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_24_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_24_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_24_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_24_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_24_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_24_BYTE_OFFSET 13'h0af8
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_25_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_25_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_25_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_25_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_25_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_25_BYTE_OFFSET 13'h0afc
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_26_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_26_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_26_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_26_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_26_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_26_BYTE_OFFSET 13'h0b00
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_27_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_27_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_27_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_27_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_27_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_27_BYTE_OFFSET 13'h0b04
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_28_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_28_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_28_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_28_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_28_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_28_BYTE_OFFSET 13'h0b08
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_29_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_29_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_29_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_29_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_29_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_29_BYTE_OFFSET 13'h0b0c
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_30_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_30_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_30_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_30_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_30_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_30_BYTE_OFFSET 13'h0b10
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_31_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_31_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_31_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_31_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_31_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_31_BYTE_OFFSET 13'h0b14
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_32_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_32_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_32_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_32_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_32_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_32_BYTE_OFFSET 13'h0b18
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_33_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_33_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_33_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_33_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_33_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_33_BYTE_OFFSET 13'h0b1c
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_34_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_34_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_34_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_34_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_34_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_34_BYTE_OFFSET 13'h0b20
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_35_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_35_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_35_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_35_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_35_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_35_BYTE_OFFSET 13'h0b24
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_36_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_36_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_36_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_36_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_36_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_36_BYTE_OFFSET 13'h0b28
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_37_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_37_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_37_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_37_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_37_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_37_BYTE_OFFSET 13'h0b2c
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_38_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_38_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_38_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_38_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_38_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_38_BYTE_OFFSET 13'h0b30
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_39_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_39_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_39_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_39_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_39_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_39_BYTE_OFFSET 13'h0b34
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_40_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_40_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_40_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_40_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_40_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_40_BYTE_OFFSET 13'h0b38
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_41_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_41_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_41_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_41_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_41_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_41_BYTE_OFFSET 13'h0b3c
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_42_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_42_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_42_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_42_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_42_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_42_BYTE_OFFSET 13'h0b40
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_43_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_43_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_43_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_43_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_43_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_43_BYTE_OFFSET 13'h0b44
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_44_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_44_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_44_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_44_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_44_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_44_BYTE_OFFSET 13'h0b48
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_45_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_45_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_45_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_45_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_45_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_45_BYTE_OFFSET 13'h0b4c
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_46_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_46_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_46_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_46_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_46_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_46_BYTE_OFFSET 13'h0b50
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_47_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_47_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_47_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_47_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_47_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_47_BYTE_OFFSET 13'h0b54
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_48_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_48_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_48_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_48_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_48_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_48_BYTE_OFFSET 13'h0b58
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_49_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_49_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_49_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_49_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_49_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_49_BYTE_OFFSET 13'h0b5c
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_50_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_50_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_50_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_50_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_50_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_50_BYTE_OFFSET 13'h0b60
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_51_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_51_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_51_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_51_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_51_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_51_BYTE_OFFSET 13'h0b64
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_52_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_52_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_52_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_52_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_52_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_52_BYTE_OFFSET 13'h0b68
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_53_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_53_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_53_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_53_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_53_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_53_BYTE_OFFSET 13'h0b6c
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_54_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_54_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_54_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_54_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_54_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_54_BYTE_OFFSET 13'h0b70
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_55_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_55_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_55_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_55_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_55_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_55_BYTE_OFFSET 13'h0b74
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_56_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_56_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_56_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_56_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_56_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_56_BYTE_OFFSET 13'h0b78
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_57_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_57_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_57_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_57_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_57_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_57_BYTE_OFFSET 13'h0b7c
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_58_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_58_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_58_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_58_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_58_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_58_BYTE_OFFSET 13'h0b80
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_59_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_59_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_59_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_59_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_59_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_59_BYTE_OFFSET 13'h0b84
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_60_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_60_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_60_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_60_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_60_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_60_BYTE_OFFSET 13'h0b88
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_61_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_61_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_61_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_61_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_61_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_61_BYTE_OFFSET 13'h0b8c
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_62_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_62_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_62_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_62_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_62_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_62_BYTE_OFFSET 13'h0b90
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_63_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_63_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_63_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_63_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_63_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_63_BYTE_OFFSET 13'h0b94
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_64_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_64_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_64_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_64_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_64_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_64_BYTE_OFFSET 13'h0b98
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_65_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_65_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_65_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_65_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_65_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_65_BYTE_OFFSET 13'h0b9c
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_66_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_66_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_66_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_66_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_66_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_66_BYTE_OFFSET 13'h0ba0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_67_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_67_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_67_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_67_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_67_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_67_BYTE_OFFSET 13'h0ba4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_68_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_68_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_68_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_68_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_68_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_68_BYTE_OFFSET 13'h0ba8
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_69_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_69_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_69_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_69_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_69_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_69_BYTE_OFFSET 13'h0bac
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_70_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_70_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_70_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_70_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_70_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_70_BYTE_OFFSET 13'h0bb0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_71_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_71_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_71_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_71_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_71_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_71_BYTE_OFFSET 13'h0bb4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_72_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_72_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_72_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_72_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_72_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_72_BYTE_OFFSET 13'h0bb8
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_73_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_73_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_73_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_73_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_73_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_73_BYTE_OFFSET 13'h0bbc
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_74_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_74_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_74_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_74_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_74_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_74_BYTE_OFFSET 13'h0bc0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_75_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_75_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_75_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_75_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_75_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_75_BYTE_OFFSET 13'h0bc4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_76_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_76_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_76_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_76_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_76_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_76_BYTE_OFFSET 13'h0bc8
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_77_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_77_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_77_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_77_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_77_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_77_BYTE_OFFSET 13'h0bcc
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_78_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_78_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_78_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_78_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_78_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_78_BYTE_OFFSET 13'h0bd0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_79_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_79_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_79_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_79_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_79_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_79_BYTE_OFFSET 13'h0bd4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_80_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_80_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_80_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_80_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_80_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_80_BYTE_OFFSET 13'h0bd8
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_81_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_81_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_81_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_81_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_81_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_81_BYTE_OFFSET 13'h0bdc
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_82_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_82_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_82_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_82_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_82_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_82_BYTE_OFFSET 13'h0be0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_83_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_83_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_83_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_83_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_83_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_83_BYTE_OFFSET 13'h0be4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_84_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_84_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_84_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_84_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_84_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_84_BYTE_OFFSET 13'h0be8
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_85_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_85_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_85_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_85_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_85_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_85_BYTE_OFFSET 13'h0bec
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_86_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_86_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_86_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_86_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_86_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_86_BYTE_OFFSET 13'h0bf0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_87_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_87_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_87_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_87_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_87_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_87_BYTE_OFFSET 13'h0bf4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_88_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_88_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_88_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_88_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_88_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_88_BYTE_OFFSET 13'h0bf8
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_89_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_89_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_89_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_89_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_89_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_89_BYTE_OFFSET 13'h0bfc
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_90_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_90_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_90_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_90_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_90_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_90_BYTE_OFFSET 13'h0c00
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_91_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_91_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_91_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_91_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_91_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_91_BYTE_OFFSET 13'h0c04
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_92_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_92_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_92_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_92_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_92_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_92_BYTE_OFFSET 13'h0c08
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_93_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_93_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_93_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_93_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_93_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_93_BYTE_OFFSET 13'h0c0c
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_94_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_94_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_94_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_94_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_94_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_94_BYTE_OFFSET 13'h0c10
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_95_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_95_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_95_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_95_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_95_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_95_BYTE_OFFSET 13'h0c14
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_96_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_96_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_96_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_96_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_96_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_96_BYTE_OFFSET 13'h0c18
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_97_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_97_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_97_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_97_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_97_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_97_BYTE_OFFSET 13'h0c1c
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_98_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_98_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_98_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_98_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_98_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_98_BYTE_OFFSET 13'h0c20
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_99_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_99_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_99_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_99_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_99_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_99_BYTE_OFFSET 13'h0c24
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_100_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_100_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_100_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_100_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_100_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_100_BYTE_OFFSET 13'h0c28
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_101_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_101_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_101_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_101_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_101_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_101_BYTE_OFFSET 13'h0c2c
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_102_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_102_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_102_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_102_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_102_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_102_BYTE_OFFSET 13'h0c30
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_103_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_103_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_103_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_103_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_103_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_103_BYTE_OFFSET 13'h0c34
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_104_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_104_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_104_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_104_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_104_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_104_BYTE_OFFSET 13'h0c38
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_105_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_105_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_105_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_105_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_105_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_105_BYTE_OFFSET 13'h0c3c
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_106_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_106_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_106_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_106_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_106_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_106_BYTE_OFFSET 13'h0c40
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_107_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_107_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_107_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_107_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_107_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_107_BYTE_OFFSET 13'h0c44
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_108_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_108_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_108_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_108_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_108_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_108_BYTE_OFFSET 13'h0c48
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_109_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_109_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_109_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_109_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_109_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_109_BYTE_OFFSET 13'h0c4c
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_110_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_110_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_110_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_110_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_110_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_110_BYTE_OFFSET 13'h0c50
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_111_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_111_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_111_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_111_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_111_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_111_BYTE_OFFSET 13'h0c54
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_112_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_112_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_112_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_112_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_112_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_112_BYTE_OFFSET 13'h0c58
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_113_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_113_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_113_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_113_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_113_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_113_BYTE_OFFSET 13'h0c5c
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_114_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_114_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_114_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_114_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_114_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_114_BYTE_OFFSET 13'h0c60
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_115_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_115_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_115_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_115_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_115_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_115_BYTE_OFFSET 13'h0c64
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_116_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_116_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_116_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_116_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_116_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_116_BYTE_OFFSET 13'h0c68
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_117_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_117_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_117_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_117_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_117_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_117_BYTE_OFFSET 13'h0c6c
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_118_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_118_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_118_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_118_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_118_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_118_BYTE_OFFSET 13'h0c70
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_119_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_119_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_119_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_119_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_119_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_119_BYTE_OFFSET 13'h0c74
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_120_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_120_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_120_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_120_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_120_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_120_BYTE_OFFSET 13'h0c78
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_121_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_121_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_121_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_121_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_121_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_121_BYTE_OFFSET 13'h0c7c
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_122_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_122_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_122_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_122_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_122_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_122_BYTE_OFFSET 13'h0c80
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_123_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_123_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_123_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_123_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_123_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_123_BYTE_OFFSET 13'h0c84
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_124_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_124_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_124_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_124_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_124_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_124_BYTE_OFFSET 13'h0c88
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_125_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_125_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_125_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_125_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_125_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_125_BYTE_OFFSET 13'h0c8c
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_126_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_126_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_126_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_126_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_126_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_126_BYTE_OFFSET 13'h0c90
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_127_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_127_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_127_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_127_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_127_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_127_BYTE_OFFSET 13'h0c94
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_128_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_128_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_128_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_128_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_128_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_128_BYTE_OFFSET 13'h0c98
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_129_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_129_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_129_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_129_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_129_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_129_BYTE_OFFSET 13'h0c9c
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_130_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_130_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_130_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_130_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_130_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_130_BYTE_OFFSET 13'h0ca0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_131_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_131_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_131_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_131_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_131_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_131_BYTE_OFFSET 13'h0ca4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_132_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_132_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_132_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_132_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_132_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_132_BYTE_OFFSET 13'h0ca8
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_133_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_133_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_133_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_133_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_133_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_133_BYTE_OFFSET 13'h0cac
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_134_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_134_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_134_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_134_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_134_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_134_BYTE_OFFSET 13'h0cb0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_135_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_135_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_135_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_135_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_135_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_135_BYTE_OFFSET 13'h0cb4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_136_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_136_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_136_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_136_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_136_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_136_BYTE_OFFSET 13'h0cb8
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_137_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_137_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_137_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_137_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_137_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_137_BYTE_OFFSET 13'h0cbc
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_138_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_138_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_138_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_138_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_138_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_138_BYTE_OFFSET 13'h0cc0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_139_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_139_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_139_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_139_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_139_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_139_BYTE_OFFSET 13'h0cc4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_140_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_140_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_140_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_140_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_140_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_140_BYTE_OFFSET 13'h0cc8
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_141_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_141_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_141_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_141_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_141_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_141_BYTE_OFFSET 13'h0ccc
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_142_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_142_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_142_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_142_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_142_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_142_BYTE_OFFSET 13'h0cd0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_143_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_143_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_143_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_143_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_143_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_143_BYTE_OFFSET 13'h0cd4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_144_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_144_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_144_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_144_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_144_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_144_BYTE_OFFSET 13'h0cd8
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_145_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_145_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_145_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_145_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_145_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_145_BYTE_OFFSET 13'h0cdc
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_146_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_146_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_146_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_146_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_146_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_146_BYTE_OFFSET 13'h0ce0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_147_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_147_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_147_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_147_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_147_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_147_BYTE_OFFSET 13'h0ce4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_148_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_148_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_148_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_148_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_148_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_148_BYTE_OFFSET 13'h0ce8
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_149_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_149_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_149_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_149_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_149_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_149_BYTE_OFFSET 13'h0cec
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_150_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_150_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_150_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_150_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_150_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_150_BYTE_OFFSET 13'h0cf0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_151_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_151_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_151_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_151_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_151_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_151_BYTE_OFFSET 13'h0cf4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_152_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_152_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_152_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_152_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_152_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_152_BYTE_OFFSET 13'h0cf8
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_153_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_153_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_153_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_153_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_153_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_153_BYTE_OFFSET 13'h0cfc
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_154_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_154_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_154_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_154_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_154_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_154_BYTE_OFFSET 13'h0d00
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_155_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_155_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_155_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_155_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_155_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_155_BYTE_OFFSET 13'h0d04
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_156_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_156_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_156_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_156_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_156_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_156_BYTE_OFFSET 13'h0d08
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_157_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_157_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_157_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_157_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_157_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_157_BYTE_OFFSET 13'h0d0c
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_158_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_158_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_158_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_158_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_158_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_158_BYTE_OFFSET 13'h0d10
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_159_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_159_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_159_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_159_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_159_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_159_BYTE_OFFSET 13'h0d14
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_160_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_160_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_160_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_160_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_160_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_160_BYTE_OFFSET 13'h0d18
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_161_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_161_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_161_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_161_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_161_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_161_BYTE_OFFSET 13'h0d1c
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_162_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_162_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_162_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_162_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_162_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_162_BYTE_OFFSET 13'h0d20
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_163_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_163_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_163_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_163_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_163_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_163_BYTE_OFFSET 13'h0d24
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_164_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_164_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_164_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_164_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_164_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_164_BYTE_OFFSET 13'h0d28
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_165_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_165_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_165_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_165_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_165_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_165_BYTE_OFFSET 13'h0d2c
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_166_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_166_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_166_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_166_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_166_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_166_BYTE_OFFSET 13'h0d30
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_167_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_167_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_167_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_167_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_167_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_167_BYTE_OFFSET 13'h0d34
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_168_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_168_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_168_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_168_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_168_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_168_BYTE_OFFSET 13'h0d38
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_169_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_169_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_169_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_169_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_169_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_169_BYTE_OFFSET 13'h0d3c
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_170_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_170_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_170_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_170_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_170_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_170_BYTE_OFFSET 13'h0d40
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_171_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_171_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_171_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_171_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_171_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_171_BYTE_OFFSET 13'h0d44
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_172_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_172_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_172_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_172_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_172_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_172_BYTE_OFFSET 13'h0d48
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_173_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_173_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_173_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_173_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_173_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_173_BYTE_OFFSET 13'h0d4c
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_174_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_174_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_174_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_174_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_174_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_174_BYTE_OFFSET 13'h0d50
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_175_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_175_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_175_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_175_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_175_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_175_BYTE_OFFSET 13'h0d54
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_176_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_176_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_176_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_176_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_176_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_176_BYTE_OFFSET 13'h0d58
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_177_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_177_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_177_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_177_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_177_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_177_BYTE_OFFSET 13'h0d5c
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_178_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_178_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_178_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_178_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_178_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_178_BYTE_OFFSET 13'h0d60
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_179_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_179_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_179_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_179_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_179_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_179_BYTE_OFFSET 13'h0d64
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_180_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_180_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_180_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_180_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_180_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_180_BYTE_OFFSET 13'h0d68
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_181_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_181_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_181_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_181_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_181_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_181_BYTE_OFFSET 13'h0d6c
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_182_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_182_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_182_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_182_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_182_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_182_BYTE_OFFSET 13'h0d70
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_183_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_183_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_183_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_183_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_183_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_183_BYTE_OFFSET 13'h0d74
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_184_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_184_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_184_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_184_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_184_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_184_BYTE_OFFSET 13'h0d78
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_185_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_185_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_185_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_185_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_185_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_185_BYTE_OFFSET 13'h0d7c
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_186_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_186_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_186_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_186_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_186_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_186_BYTE_OFFSET 13'h0d80
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_187_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_187_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_187_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_187_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_187_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_187_BYTE_OFFSET 13'h0d84
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_188_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_188_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_188_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_188_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_188_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_188_BYTE_OFFSET 13'h0d88
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_189_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_189_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_189_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_189_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_189_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_189_BYTE_OFFSET 13'h0d8c
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_190_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_190_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_190_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_190_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_190_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_190_BYTE_OFFSET 13'h0d90
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_191_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_191_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_191_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_191_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_191_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_191_BYTE_OFFSET 13'h0d94
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_192_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_192_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_192_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_192_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_192_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_192_BYTE_OFFSET 13'h0d98
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_193_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_193_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_193_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_193_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_193_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_193_BYTE_OFFSET 13'h0d9c
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_194_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_194_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_194_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_194_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_194_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_194_BYTE_OFFSET 13'h0da0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_195_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_195_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_195_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_195_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_195_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_195_BYTE_OFFSET 13'h0da4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_196_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_196_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_196_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_196_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_196_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_196_BYTE_OFFSET 13'h0da8
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_197_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_197_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_197_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_197_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_197_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_197_BYTE_OFFSET 13'h0dac
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_198_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_198_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_198_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_198_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_198_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_198_BYTE_OFFSET 13'h0db0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_199_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_199_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_199_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_199_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_199_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_199_BYTE_OFFSET 13'h0db4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_200_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_200_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_200_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_200_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_200_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_200_BYTE_OFFSET 13'h0db8
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_201_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_201_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_201_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_201_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_201_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_201_BYTE_OFFSET 13'h0dbc
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_202_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_202_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_202_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_202_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_202_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_202_BYTE_OFFSET 13'h0dc0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_203_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_203_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_203_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_203_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_203_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_203_BYTE_OFFSET 13'h0dc4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_204_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_204_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_204_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_204_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_204_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_204_BYTE_OFFSET 13'h0dc8
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_205_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_205_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_205_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_205_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_205_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_205_BYTE_OFFSET 13'h0dcc
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_206_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_206_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_206_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_206_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_206_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_206_BYTE_OFFSET 13'h0dd0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_207_FINAL_CWORD_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_207_FINAL_CWORD_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_207_FINAL_CWORD_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_207_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_207_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_CODEWRD_OUT_BIT_207_BYTE_OFFSET 13'h0dd4
`define LDPC_CSR_LDPC_DEC_PASS_FAIL_PASS_FAIL_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_PASS_FAIL_PASS_FAIL_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_PASS_FAIL_PASS_FAIL_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_PASS_FAIL_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_PASS_FAIL_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_PASS_FAIL_BYTE_OFFSET 13'h0dd8
`define LDPC_CSR_LDPC_DEC_TB_PASS_FAIL_DECODER_TB_PASS_FAIL_DECODER_BIT_BIT_WIDTH 1
`define LDPC_CSR_LDPC_DEC_TB_PASS_FAIL_DECODER_TB_PASS_FAIL_DECODER_BIT_BIT_MASK 1'h1
`define LDPC_CSR_LDPC_DEC_TB_PASS_FAIL_DECODER_TB_PASS_FAIL_DECODER_BIT_BIT_OFFSET 0
`define LDPC_CSR_LDPC_DEC_TB_PASS_FAIL_DECODER_BYTE_WIDTH 4
`define LDPC_CSR_LDPC_DEC_TB_PASS_FAIL_DECODER_BYTE_SIZE 4
`define LDPC_CSR_LDPC_DEC_TB_PASS_FAIL_DECODER_BYTE_OFFSET 13'h0ddc
`endif
