wire o_LDPC_ENC_MSG_IN_0_msg_in;
wire o_LDPC_ENC_MSG_IN_1_msg_in;
wire o_LDPC_ENC_MSG_IN_2_msg_in;
wire o_LDPC_ENC_MSG_IN_3_msg_in;
wire o_LDPC_ENC_MSG_IN_4_msg_in;
wire o_LDPC_ENC_MSG_IN_5_msg_in;
wire o_LDPC_ENC_MSG_IN_6_msg_in;
wire o_LDPC_ENC_MSG_IN_7_msg_in;
wire o_LDPC_ENC_MSG_IN_8_msg_in;
wire o_LDPC_ENC_MSG_IN_9_msg_in;
wire o_LDPC_ENC_MSG_IN_10_msg_in;
wire o_LDPC_ENC_MSG_IN_11_msg_in;
wire o_LDPC_ENC_MSG_IN_12_msg_in;
wire o_LDPC_ENC_MSG_IN_13_msg_in;
wire o_LDPC_ENC_MSG_IN_14_msg_in;
wire o_LDPC_ENC_MSG_IN_15_msg_in;
wire o_LDPC_ENC_MSG_IN_16_msg_in;
wire o_LDPC_ENC_MSG_IN_17_msg_in;
wire o_LDPC_ENC_MSG_IN_18_msg_in;
wire o_LDPC_ENC_MSG_IN_19_msg_in;
wire o_LDPC_ENC_MSG_IN_20_msg_in;
wire o_LDPC_ENC_MSG_IN_21_msg_in;
wire o_LDPC_ENC_MSG_IN_22_msg_in;
wire o_LDPC_ENC_MSG_IN_23_msg_in;
wire o_LDPC_ENC_MSG_IN_24_msg_in;
wire o_LDPC_ENC_MSG_IN_25_msg_in;
wire o_LDPC_ENC_MSG_IN_26_msg_in;
wire o_LDPC_ENC_MSG_IN_27_msg_in;
wire o_LDPC_ENC_MSG_IN_28_msg_in;
wire o_LDPC_ENC_MSG_IN_29_msg_in;
wire o_LDPC_ENC_MSG_IN_30_msg_in;
wire o_LDPC_ENC_MSG_IN_31_msg_in;
wire o_LDPC_ENC_MSG_IN_32_msg_in;
wire o_LDPC_ENC_MSG_IN_33_msg_in;
wire o_LDPC_ENC_MSG_IN_34_msg_in;
wire o_LDPC_ENC_MSG_IN_35_msg_in;
wire o_LDPC_ENC_MSG_IN_36_msg_in;
wire o_LDPC_ENC_MSG_IN_37_msg_in;
wire o_LDPC_ENC_MSG_IN_38_msg_in;
wire o_LDPC_ENC_MSG_IN_39_msg_in;
wire i_LDPC_ENC_CODEWRD_0_enc_codeword;
wire i_LDPC_ENC_CODEWRD_1_enc_codeword;
wire i_LDPC_ENC_CODEWRD_2_enc_codeword;
wire i_LDPC_ENC_CODEWRD_3_enc_codeword;
wire i_LDPC_ENC_CODEWRD_4_enc_codeword;
wire i_LDPC_ENC_CODEWRD_5_enc_codeword;
wire i_LDPC_ENC_CODEWRD_6_enc_codeword;
wire i_LDPC_ENC_CODEWRD_7_enc_codeword;
wire i_LDPC_ENC_CODEWRD_8_enc_codeword;
wire i_LDPC_ENC_CODEWRD_9_enc_codeword;
wire i_LDPC_ENC_CODEWRD_10_enc_codeword;
wire i_LDPC_ENC_CODEWRD_11_enc_codeword;
wire i_LDPC_ENC_CODEWRD_12_enc_codeword;
wire i_LDPC_ENC_CODEWRD_13_enc_codeword;
wire i_LDPC_ENC_CODEWRD_14_enc_codeword;
wire i_LDPC_ENC_CODEWRD_15_enc_codeword;
wire i_LDPC_ENC_CODEWRD_16_enc_codeword;
wire i_LDPC_ENC_CODEWRD_17_enc_codeword;
wire i_LDPC_ENC_CODEWRD_18_enc_codeword;
wire i_LDPC_ENC_CODEWRD_19_enc_codeword;
wire i_LDPC_ENC_CODEWRD_20_enc_codeword;
wire i_LDPC_ENC_CODEWRD_21_enc_codeword;
wire i_LDPC_ENC_CODEWRD_22_enc_codeword;
wire i_LDPC_ENC_CODEWRD_23_enc_codeword;
wire i_LDPC_ENC_CODEWRD_24_enc_codeword;
wire i_LDPC_ENC_CODEWRD_25_enc_codeword;
wire i_LDPC_ENC_CODEWRD_26_enc_codeword;
wire i_LDPC_ENC_CODEWRD_27_enc_codeword;
wire i_LDPC_ENC_CODEWRD_28_enc_codeword;
wire i_LDPC_ENC_CODEWRD_29_enc_codeword;
wire i_LDPC_ENC_CODEWRD_30_enc_codeword;
wire i_LDPC_ENC_CODEWRD_31_enc_codeword;
wire i_LDPC_ENC_CODEWRD_32_enc_codeword;
wire i_LDPC_ENC_CODEWRD_33_enc_codeword;
wire i_LDPC_ENC_CODEWRD_34_enc_codeword;
wire i_LDPC_ENC_CODEWRD_35_enc_codeword;
wire i_LDPC_ENC_CODEWRD_36_enc_codeword;
wire i_LDPC_ENC_CODEWRD_37_enc_codeword;
wire i_LDPC_ENC_CODEWRD_38_enc_codeword;
wire i_LDPC_ENC_CODEWRD_39_enc_codeword;
wire i_LDPC_ENC_CODEWRD_40_enc_codeword;
wire i_LDPC_ENC_CODEWRD_41_enc_codeword;
wire i_LDPC_ENC_CODEWRD_42_enc_codeword;
wire i_LDPC_ENC_CODEWRD_43_enc_codeword;
wire i_LDPC_ENC_CODEWRD_44_enc_codeword;
wire i_LDPC_ENC_CODEWRD_45_enc_codeword;
wire i_LDPC_ENC_CODEWRD_46_enc_codeword;
wire i_LDPC_ENC_CODEWRD_47_enc_codeword;
wire i_LDPC_ENC_CODEWRD_48_enc_codeword;
wire i_LDPC_ENC_CODEWRD_49_enc_codeword;
wire i_LDPC_ENC_CODEWRD_50_enc_codeword;
wire i_LDPC_ENC_CODEWRD_51_enc_codeword;
wire i_LDPC_ENC_CODEWRD_52_enc_codeword;
wire i_LDPC_ENC_CODEWRD_53_enc_codeword;
wire i_LDPC_ENC_CODEWRD_54_enc_codeword;
wire i_LDPC_ENC_CODEWRD_55_enc_codeword;
wire i_LDPC_ENC_CODEWRD_56_enc_codeword;
wire i_LDPC_ENC_CODEWRD_57_enc_codeword;
wire i_LDPC_ENC_CODEWRD_58_enc_codeword;
wire i_LDPC_ENC_CODEWRD_59_enc_codeword;
wire i_LDPC_ENC_CODEWRD_60_enc_codeword;
wire i_LDPC_ENC_CODEWRD_61_enc_codeword;
wire i_LDPC_ENC_CODEWRD_62_enc_codeword;
wire i_LDPC_ENC_CODEWRD_63_enc_codeword;
wire i_LDPC_ENC_CODEWRD_64_enc_codeword;
wire i_LDPC_ENC_CODEWRD_65_enc_codeword;
wire i_LDPC_ENC_CODEWRD_66_enc_codeword;
wire i_LDPC_ENC_CODEWRD_67_enc_codeword;
wire i_LDPC_ENC_CODEWRD_68_enc_codeword;
wire i_LDPC_ENC_CODEWRD_69_enc_codeword;
wire i_LDPC_ENC_CODEWRD_70_enc_codeword;
wire i_LDPC_ENC_CODEWRD_71_enc_codeword;
wire i_LDPC_ENC_CODEWRD_72_enc_codeword;
wire i_LDPC_ENC_CODEWRD_73_enc_codeword;
wire i_LDPC_ENC_CODEWRD_74_enc_codeword;
wire i_LDPC_ENC_CODEWRD_75_enc_codeword;
wire i_LDPC_ENC_CODEWRD_76_enc_codeword;
wire i_LDPC_ENC_CODEWRD_77_enc_codeword;
wire i_LDPC_ENC_CODEWRD_78_enc_codeword;
wire i_LDPC_ENC_CODEWRD_79_enc_codeword;
wire i_LDPC_ENC_CODEWRD_80_enc_codeword;
wire i_LDPC_ENC_CODEWRD_81_enc_codeword;
wire i_LDPC_ENC_CODEWRD_82_enc_codeword;
wire i_LDPC_ENC_CODEWRD_83_enc_codeword;
wire i_LDPC_ENC_CODEWRD_84_enc_codeword;
wire i_LDPC_ENC_CODEWRD_85_enc_codeword;
wire i_LDPC_ENC_CODEWRD_86_enc_codeword;
wire i_LDPC_ENC_CODEWRD_87_enc_codeword;
wire i_LDPC_ENC_CODEWRD_88_enc_codeword;
wire i_LDPC_ENC_CODEWRD_89_enc_codeword;
wire i_LDPC_ENC_CODEWRD_90_enc_codeword;
wire i_LDPC_ENC_CODEWRD_91_enc_codeword;
wire i_LDPC_ENC_CODEWRD_92_enc_codeword;
wire i_LDPC_ENC_CODEWRD_93_enc_codeword;
wire i_LDPC_ENC_CODEWRD_94_enc_codeword;
wire i_LDPC_ENC_CODEWRD_95_enc_codeword;
wire i_LDPC_ENC_CODEWRD_96_enc_codeword;
wire i_LDPC_ENC_CODEWRD_97_enc_codeword;
wire i_LDPC_ENC_CODEWRD_98_enc_codeword;
wire i_LDPC_ENC_CODEWRD_99_enc_codeword;
wire i_LDPC_ENC_CODEWRD_100_enc_codeword;
wire i_LDPC_ENC_CODEWRD_101_enc_codeword;
wire i_LDPC_ENC_CODEWRD_102_enc_codeword;
wire i_LDPC_ENC_CODEWRD_103_enc_codeword;
wire i_LDPC_ENC_CODEWRD_104_enc_codeword;
wire i_LDPC_ENC_CODEWRD_105_enc_codeword;
wire i_LDPC_ENC_CODEWRD_106_enc_codeword;
wire i_LDPC_ENC_CODEWRD_107_enc_codeword;
wire i_LDPC_ENC_CODEWRD_108_enc_codeword;
wire i_LDPC_ENC_CODEWRD_109_enc_codeword;
wire i_LDPC_ENC_CODEWRD_110_enc_codeword;
wire i_LDPC_ENC_CODEWRD_111_enc_codeword;
wire i_LDPC_ENC_CODEWRD_112_enc_codeword;
wire i_LDPC_ENC_CODEWRD_113_enc_codeword;
wire i_LDPC_ENC_CODEWRD_114_enc_codeword;
wire i_LDPC_ENC_CODEWRD_115_enc_codeword;
wire i_LDPC_ENC_CODEWRD_116_enc_codeword;
wire i_LDPC_ENC_CODEWRD_117_enc_codeword;
wire i_LDPC_ENC_CODEWRD_118_enc_codeword;
wire i_LDPC_ENC_CODEWRD_119_enc_codeword;
wire i_LDPC_ENC_CODEWRD_120_enc_codeword;
wire i_LDPC_ENC_CODEWRD_121_enc_codeword;
wire i_LDPC_ENC_CODEWRD_122_enc_codeword;
wire i_LDPC_ENC_CODEWRD_123_enc_codeword;
wire i_LDPC_ENC_CODEWRD_124_enc_codeword;
wire i_LDPC_ENC_CODEWRD_125_enc_codeword;
wire i_LDPC_ENC_CODEWRD_126_enc_codeword;
wire i_LDPC_ENC_CODEWRD_127_enc_codeword;
wire i_LDPC_ENC_CODEWRD_128_enc_codeword;
wire i_LDPC_ENC_CODEWRD_129_enc_codeword;
wire i_LDPC_ENC_CODEWRD_130_enc_codeword;
wire i_LDPC_ENC_CODEWRD_131_enc_codeword;
wire i_LDPC_ENC_CODEWRD_132_enc_codeword;
wire i_LDPC_ENC_CODEWRD_133_enc_codeword;
wire i_LDPC_ENC_CODEWRD_134_enc_codeword;
wire i_LDPC_ENC_CODEWRD_135_enc_codeword;
wire i_LDPC_ENC_CODEWRD_136_enc_codeword;
wire i_LDPC_ENC_CODEWRD_137_enc_codeword;
wire i_LDPC_ENC_CODEWRD_138_enc_codeword;
wire i_LDPC_ENC_CODEWRD_139_enc_codeword;
wire i_LDPC_ENC_CODEWRD_140_enc_codeword;
wire i_LDPC_ENC_CODEWRD_141_enc_codeword;
wire i_LDPC_ENC_CODEWRD_142_enc_codeword;
wire i_LDPC_ENC_CODEWRD_143_enc_codeword;
wire i_LDPC_ENC_CODEWRD_144_enc_codeword;
wire i_LDPC_ENC_CODEWRD_145_enc_codeword;
wire i_LDPC_ENC_CODEWRD_146_enc_codeword;
wire i_LDPC_ENC_CODEWRD_147_enc_codeword;
wire i_LDPC_ENC_CODEWRD_148_enc_codeword;
wire i_LDPC_ENC_CODEWRD_149_enc_codeword;
wire i_LDPC_ENC_CODEWRD_150_enc_codeword;
wire i_LDPC_ENC_CODEWRD_151_enc_codeword;
wire i_LDPC_ENC_CODEWRD_152_enc_codeword;
wire i_LDPC_ENC_CODEWRD_153_enc_codeword;
wire i_LDPC_ENC_CODEWRD_154_enc_codeword;
wire i_LDPC_ENC_CODEWRD_155_enc_codeword;
wire i_LDPC_ENC_CODEWRD_156_enc_codeword;
wire i_LDPC_ENC_CODEWRD_157_enc_codeword;
wire i_LDPC_ENC_CODEWRD_158_enc_codeword;
wire i_LDPC_ENC_CODEWRD_159_enc_codeword;
wire i_LDPC_ENC_CODEWRD_160_enc_codeword;
wire i_LDPC_ENC_CODEWRD_161_enc_codeword;
wire i_LDPC_ENC_CODEWRD_162_enc_codeword;
wire i_LDPC_ENC_CODEWRD_163_enc_codeword;
wire i_LDPC_ENC_CODEWRD_164_enc_codeword;
wire i_LDPC_ENC_CODEWRD_165_enc_codeword;
wire i_LDPC_ENC_CODEWRD_166_enc_codeword;
wire i_LDPC_ENC_CODEWRD_167_enc_codeword;
wire i_LDPC_ENC_CODEWRD_168_enc_codeword;
wire i_LDPC_ENC_CODEWRD_169_enc_codeword;
wire i_LDPC_ENC_CODEWRD_170_enc_codeword;
wire i_LDPC_ENC_CODEWRD_171_enc_codeword;
wire i_LDPC_ENC_CODEWRD_172_enc_codeword;
wire i_LDPC_ENC_CODEWRD_173_enc_codeword;
wire i_LDPC_ENC_CODEWRD_174_enc_codeword;
wire i_LDPC_ENC_CODEWRD_175_enc_codeword;
wire i_LDPC_ENC_CODEWRD_176_enc_codeword;
wire i_LDPC_ENC_CODEWRD_177_enc_codeword;
wire i_LDPC_ENC_CODEWRD_178_enc_codeword;
wire i_LDPC_ENC_CODEWRD_179_enc_codeword;
wire i_LDPC_ENC_CODEWRD_180_enc_codeword;
wire i_LDPC_ENC_CODEWRD_181_enc_codeword;
wire i_LDPC_ENC_CODEWRD_182_enc_codeword;
wire i_LDPC_ENC_CODEWRD_183_enc_codeword;
wire i_LDPC_ENC_CODEWRD_184_enc_codeword;
wire i_LDPC_ENC_CODEWRD_185_enc_codeword;
wire i_LDPC_ENC_CODEWRD_186_enc_codeword;
wire i_LDPC_ENC_CODEWRD_187_enc_codeword;
wire i_LDPC_ENC_CODEWRD_188_enc_codeword;
wire i_LDPC_ENC_CODEWRD_189_enc_codeword;
wire i_LDPC_ENC_CODEWRD_190_enc_codeword;
wire i_LDPC_ENC_CODEWRD_191_enc_codeword;
wire i_LDPC_ENC_CODEWRD_192_enc_codeword;
wire i_LDPC_ENC_CODEWRD_193_enc_codeword;
wire i_LDPC_ENC_CODEWRD_194_enc_codeword;
wire i_LDPC_ENC_CODEWRD_195_enc_codeword;
wire i_LDPC_ENC_CODEWRD_196_enc_codeword;
wire i_LDPC_ENC_CODEWRD_197_enc_codeword;
wire i_LDPC_ENC_CODEWRD_198_enc_codeword;
wire i_LDPC_ENC_CODEWRD_199_enc_codeword;
wire i_LDPC_ENC_CODEWRD_200_enc_codeword;
wire i_LDPC_ENC_CODEWRD_201_enc_codeword;
wire i_LDPC_ENC_CODEWRD_202_enc_codeword;
wire i_LDPC_ENC_CODEWRD_203_enc_codeword;
wire i_LDPC_ENC_CODEWRD_204_enc_codeword;
wire i_LDPC_ENC_CODEWRD_205_enc_codeword;
wire i_LDPC_ENC_CODEWRD_206_enc_codeword;
wire i_LDPC_ENC_CODEWRD_207_enc_codeword;
wire i_LDPC_ENC_CODEWRD_VLD_enc_codeword_valid;
wire [1:0] o_LDPC_DEC_CODEWRD_0_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_1_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_2_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_3_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_4_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_5_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_6_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_7_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_8_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_9_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_10_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_11_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_12_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_13_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_14_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_15_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_16_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_17_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_18_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_19_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_20_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_21_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_22_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_23_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_24_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_25_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_26_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_27_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_28_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_29_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_30_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_31_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_32_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_33_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_34_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_35_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_36_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_37_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_38_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_39_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_40_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_41_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_42_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_43_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_44_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_45_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_46_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_47_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_48_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_49_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_50_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_51_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_52_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_53_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_54_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_55_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_56_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_57_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_58_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_59_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_60_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_61_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_62_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_63_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_64_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_65_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_66_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_67_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_68_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_69_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_70_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_71_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_72_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_73_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_74_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_75_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_76_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_77_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_78_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_79_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_80_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_81_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_82_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_83_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_84_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_85_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_86_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_87_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_88_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_89_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_90_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_91_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_92_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_93_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_94_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_95_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_96_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_97_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_98_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_99_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_100_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_101_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_102_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_103_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_104_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_105_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_106_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_107_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_108_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_109_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_110_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_111_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_112_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_113_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_114_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_115_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_116_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_117_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_118_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_119_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_120_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_121_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_122_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_123_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_124_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_125_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_126_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_127_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_128_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_129_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_130_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_131_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_132_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_133_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_134_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_135_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_136_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_137_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_138_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_139_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_140_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_141_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_142_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_143_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_144_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_145_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_146_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_147_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_148_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_149_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_150_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_151_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_152_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_153_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_154_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_155_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_156_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_157_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_158_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_159_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_160_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_161_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_162_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_163_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_164_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_165_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_166_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_167_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_168_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_169_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_170_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_171_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_172_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_173_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_174_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_175_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_176_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_177_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_178_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_179_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_180_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_181_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_182_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_183_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_184_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_185_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_186_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_187_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_188_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_189_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_190_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_191_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_192_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_193_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_194_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_195_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_196_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_197_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_198_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_199_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_200_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_201_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_202_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_203_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_204_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_205_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_206_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_207_cword_q0;
wire o_LDPC_DEC_EXPSYND_0_exp_syn;
wire o_LDPC_DEC_EXPSYND_1_exp_syn;
wire o_LDPC_DEC_EXPSYND_2_exp_syn;
wire o_LDPC_DEC_EXPSYND_3_exp_syn;
wire o_LDPC_DEC_EXPSYND_4_exp_syn;
wire o_LDPC_DEC_EXPSYND_5_exp_syn;
wire o_LDPC_DEC_EXPSYND_6_exp_syn;
wire o_LDPC_DEC_EXPSYND_7_exp_syn;
wire o_LDPC_DEC_EXPSYND_8_exp_syn;
wire o_LDPC_DEC_EXPSYND_9_exp_syn;
wire o_LDPC_DEC_EXPSYND_10_exp_syn;
wire o_LDPC_DEC_EXPSYND_11_exp_syn;
wire o_LDPC_DEC_EXPSYND_12_exp_syn;
wire o_LDPC_DEC_EXPSYND_13_exp_syn;
wire o_LDPC_DEC_EXPSYND_14_exp_syn;
wire o_LDPC_DEC_EXPSYND_15_exp_syn;
wire o_LDPC_DEC_EXPSYND_16_exp_syn;
wire o_LDPC_DEC_EXPSYND_17_exp_syn;
wire o_LDPC_DEC_EXPSYND_18_exp_syn;
wire o_LDPC_DEC_EXPSYND_19_exp_syn;
wire o_LDPC_DEC_EXPSYND_20_exp_syn;
wire o_LDPC_DEC_EXPSYND_21_exp_syn;
wire o_LDPC_DEC_EXPSYND_22_exp_syn;
wire o_LDPC_DEC_EXPSYND_23_exp_syn;
wire o_LDPC_DEC_EXPSYND_24_exp_syn;
wire o_LDPC_DEC_EXPSYND_25_exp_syn;
wire o_LDPC_DEC_EXPSYND_26_exp_syn;
wire o_LDPC_DEC_EXPSYND_27_exp_syn;
wire o_LDPC_DEC_EXPSYND_28_exp_syn;
wire o_LDPC_DEC_EXPSYND_29_exp_syn;
wire o_LDPC_DEC_EXPSYND_30_exp_syn;
wire o_LDPC_DEC_EXPSYND_31_exp_syn;
wire o_LDPC_DEC_EXPSYND_32_exp_syn;
wire o_LDPC_DEC_EXPSYND_33_exp_syn;
wire o_LDPC_DEC_EXPSYND_34_exp_syn;
wire o_LDPC_DEC_EXPSYND_35_exp_syn;
wire o_LDPC_DEC_EXPSYND_36_exp_syn;
wire o_LDPC_DEC_EXPSYND_37_exp_syn;
wire o_LDPC_DEC_EXPSYND_38_exp_syn;
wire o_LDPC_DEC_EXPSYND_39_exp_syn;
wire o_LDPC_DEC_EXPSYND_40_exp_syn;
wire o_LDPC_DEC_EXPSYND_41_exp_syn;
wire o_LDPC_DEC_EXPSYND_42_exp_syn;
wire o_LDPC_DEC_EXPSYND_43_exp_syn;
wire o_LDPC_DEC_EXPSYND_44_exp_syn;
wire o_LDPC_DEC_EXPSYND_45_exp_syn;
wire o_LDPC_DEC_EXPSYND_46_exp_syn;
wire o_LDPC_DEC_EXPSYND_47_exp_syn;
wire o_LDPC_DEC_EXPSYND_48_exp_syn;
wire o_LDPC_DEC_EXPSYND_49_exp_syn;
wire o_LDPC_DEC_EXPSYND_50_exp_syn;
wire o_LDPC_DEC_EXPSYND_51_exp_syn;
wire o_LDPC_DEC_EXPSYND_52_exp_syn;
wire o_LDPC_DEC_EXPSYND_53_exp_syn;
wire o_LDPC_DEC_EXPSYND_54_exp_syn;
wire o_LDPC_DEC_EXPSYND_55_exp_syn;
wire o_LDPC_DEC_EXPSYND_56_exp_syn;
wire o_LDPC_DEC_EXPSYND_57_exp_syn;
wire o_LDPC_DEC_EXPSYND_58_exp_syn;
wire o_LDPC_DEC_EXPSYND_59_exp_syn;
wire o_LDPC_DEC_EXPSYND_60_exp_syn;
wire o_LDPC_DEC_EXPSYND_61_exp_syn;
wire o_LDPC_DEC_EXPSYND_62_exp_syn;
wire o_LDPC_DEC_EXPSYND_63_exp_syn;
wire o_LDPC_DEC_EXPSYND_64_exp_syn;
wire o_LDPC_DEC_EXPSYND_65_exp_syn;
wire o_LDPC_DEC_EXPSYND_66_exp_syn;
wire o_LDPC_DEC_EXPSYND_67_exp_syn;
wire o_LDPC_DEC_EXPSYND_68_exp_syn;
wire o_LDPC_DEC_EXPSYND_69_exp_syn;
wire o_LDPC_DEC_EXPSYND_70_exp_syn;
wire o_LDPC_DEC_EXPSYND_71_exp_syn;
wire o_LDPC_DEC_EXPSYND_72_exp_syn;
wire o_LDPC_DEC_EXPSYND_73_exp_syn;
wire o_LDPC_DEC_EXPSYND_74_exp_syn;
wire o_LDPC_DEC_EXPSYND_75_exp_syn;
wire o_LDPC_DEC_EXPSYND_76_exp_syn;
wire o_LDPC_DEC_EXPSYND_77_exp_syn;
wire o_LDPC_DEC_EXPSYND_78_exp_syn;
wire o_LDPC_DEC_EXPSYND_79_exp_syn;
wire o_LDPC_DEC_EXPSYND_80_exp_syn;
wire o_LDPC_DEC_EXPSYND_81_exp_syn;
wire o_LDPC_DEC_EXPSYND_82_exp_syn;
wire o_LDPC_DEC_EXPSYND_83_exp_syn;
wire o_LDPC_DEC_EXPSYND_84_exp_syn;
wire o_LDPC_DEC_EXPSYND_85_exp_syn;
wire o_LDPC_DEC_EXPSYND_86_exp_syn;
wire o_LDPC_DEC_EXPSYND_87_exp_syn;
wire o_LDPC_DEC_EXPSYND_88_exp_syn;
wire o_LDPC_DEC_EXPSYND_89_exp_syn;
wire o_LDPC_DEC_EXPSYND_90_exp_syn;
wire o_LDPC_DEC_EXPSYND_91_exp_syn;
wire o_LDPC_DEC_EXPSYND_92_exp_syn;
wire o_LDPC_DEC_EXPSYND_93_exp_syn;
wire o_LDPC_DEC_EXPSYND_94_exp_syn;
wire o_LDPC_DEC_EXPSYND_95_exp_syn;
wire o_LDPC_DEC_EXPSYND_96_exp_syn;
wire o_LDPC_DEC_EXPSYND_97_exp_syn;
wire o_LDPC_DEC_EXPSYND_98_exp_syn;
wire o_LDPC_DEC_EXPSYND_99_exp_syn;
wire o_LDPC_DEC_EXPSYND_100_exp_syn;
wire o_LDPC_DEC_EXPSYND_101_exp_syn;
wire o_LDPC_DEC_EXPSYND_102_exp_syn;
wire o_LDPC_DEC_EXPSYND_103_exp_syn;
wire o_LDPC_DEC_EXPSYND_104_exp_syn;
wire o_LDPC_DEC_EXPSYND_105_exp_syn;
wire o_LDPC_DEC_EXPSYND_106_exp_syn;
wire o_LDPC_DEC_EXPSYND_107_exp_syn;
wire o_LDPC_DEC_EXPSYND_108_exp_syn;
wire o_LDPC_DEC_EXPSYND_109_exp_syn;
wire o_LDPC_DEC_EXPSYND_110_exp_syn;
wire o_LDPC_DEC_EXPSYND_111_exp_syn;
wire o_LDPC_DEC_EXPSYND_112_exp_syn;
wire o_LDPC_DEC_EXPSYND_113_exp_syn;
wire o_LDPC_DEC_EXPSYND_114_exp_syn;
wire o_LDPC_DEC_EXPSYND_115_exp_syn;
wire o_LDPC_DEC_EXPSYND_116_exp_syn;
wire o_LDPC_DEC_EXPSYND_117_exp_syn;
wire o_LDPC_DEC_EXPSYND_118_exp_syn;
wire o_LDPC_DEC_EXPSYND_119_exp_syn;
wire o_LDPC_DEC_EXPSYND_120_exp_syn;
wire o_LDPC_DEC_EXPSYND_121_exp_syn;
wire o_LDPC_DEC_EXPSYND_122_exp_syn;
wire o_LDPC_DEC_EXPSYND_123_exp_syn;
wire o_LDPC_DEC_EXPSYND_124_exp_syn;
wire o_LDPC_DEC_EXPSYND_125_exp_syn;
wire o_LDPC_DEC_EXPSYND_126_exp_syn;
wire o_LDPC_DEC_EXPSYND_127_exp_syn;
wire o_LDPC_DEC_EXPSYND_128_exp_syn;
wire o_LDPC_DEC_EXPSYND_129_exp_syn;
wire o_LDPC_DEC_EXPSYND_130_exp_syn;
wire o_LDPC_DEC_EXPSYND_131_exp_syn;
wire o_LDPC_DEC_EXPSYND_132_exp_syn;
wire o_LDPC_DEC_EXPSYND_133_exp_syn;
wire o_LDPC_DEC_EXPSYND_134_exp_syn;
wire o_LDPC_DEC_EXPSYND_135_exp_syn;
wire o_LDPC_DEC_EXPSYND_136_exp_syn;
wire o_LDPC_DEC_EXPSYND_137_exp_syn;
wire o_LDPC_DEC_EXPSYND_138_exp_syn;
wire o_LDPC_DEC_EXPSYND_139_exp_syn;
wire o_LDPC_DEC_EXPSYND_140_exp_syn;
wire o_LDPC_DEC_EXPSYND_141_exp_syn;
wire o_LDPC_DEC_EXPSYND_142_exp_syn;
wire o_LDPC_DEC_EXPSYND_143_exp_syn;
wire o_LDPC_DEC_EXPSYND_144_exp_syn;
wire o_LDPC_DEC_EXPSYND_145_exp_syn;
wire o_LDPC_DEC_EXPSYND_146_exp_syn;
wire o_LDPC_DEC_EXPSYND_147_exp_syn;
wire o_LDPC_DEC_EXPSYND_148_exp_syn;
wire o_LDPC_DEC_EXPSYND_149_exp_syn;
wire o_LDPC_DEC_EXPSYND_150_exp_syn;
wire o_LDPC_DEC_EXPSYND_151_exp_syn;
wire o_LDPC_DEC_EXPSYND_152_exp_syn;
wire o_LDPC_DEC_EXPSYND_153_exp_syn;
wire o_LDPC_DEC_EXPSYND_154_exp_syn;
wire o_LDPC_DEC_EXPSYND_155_exp_syn;
wire o_LDPC_DEC_EXPSYND_156_exp_syn;
wire o_LDPC_DEC_EXPSYND_157_exp_syn;
wire o_LDPC_DEC_EXPSYND_158_exp_syn;
wire o_LDPC_DEC_EXPSYND_159_exp_syn;
wire o_LDPC_DEC_EXPSYND_160_exp_syn;
wire o_LDPC_DEC_EXPSYND_161_exp_syn;
wire o_LDPC_DEC_EXPSYND_162_exp_syn;
wire o_LDPC_DEC_EXPSYND_163_exp_syn;
wire o_LDPC_DEC_EXPSYND_164_exp_syn;
wire o_LDPC_DEC_EXPSYND_165_exp_syn;
wire o_LDPC_DEC_EXPSYND_166_exp_syn;
wire o_LDPC_DEC_EXPSYND_167_exp_syn;
wire [31:0] o_LDPC_DEC_PROBABILITY_perc_probability;
wire [31:0] o_LDPC_DEC_HamDist_loop_max_HamDist_loop_max;
wire [31:0] o_LDPC_DEC_HamDist_loop_percentage_HamDist_loop_percentage;
wire [31:0] o_LDPC_DEC_HamDist_iir1_HamDist_iir1;
wire [31:0] o_LDPC_DEC_HamDist_iir2_NOT_USED_HamDist_iir2;
wire [31:0] o_LDPC_DEC_HamDist_iir3_NOT_USED_HamDist_iir3;
wire i_LDPC_DEC_converged_valid_NOT_USED_convered_valid;
wire i_LDPC_DEC_valid_NOT_USED_dec_valid;
wire i_LDPC_DEC_valid_codeword_NOT_USED_dec_valid_cword;
wire o_LDPC_DEC_start_start;
wire i_LDPC_DEC_converged_valid_convered_vld;
wire i_LDPC_DEC_converged_status_convered_stat;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_0_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_1_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_2_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_3_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_4_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_5_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_6_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_7_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_8_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_9_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_10_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_11_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_12_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_13_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_14_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_15_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_16_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_17_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_18_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_19_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_20_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_21_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_22_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_23_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_24_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_25_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_26_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_27_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_28_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_29_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_30_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_31_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_32_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_33_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_34_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_35_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_36_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_37_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_38_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_39_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_40_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_41_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_42_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_43_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_44_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_45_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_46_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_47_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_48_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_49_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_50_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_51_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_52_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_53_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_54_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_55_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_56_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_57_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_58_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_59_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_60_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_61_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_62_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_63_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_64_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_65_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_66_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_67_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_68_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_69_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_70_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_71_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_72_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_73_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_74_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_75_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_76_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_77_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_78_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_79_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_80_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_81_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_82_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_83_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_84_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_85_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_86_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_87_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_88_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_89_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_90_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_91_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_92_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_93_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_94_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_95_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_96_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_97_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_98_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_99_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_100_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_101_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_102_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_103_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_104_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_105_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_106_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_107_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_108_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_109_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_110_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_111_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_112_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_113_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_114_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_115_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_116_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_117_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_118_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_119_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_120_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_121_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_122_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_123_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_124_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_125_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_126_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_127_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_128_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_129_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_130_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_131_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_132_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_133_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_134_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_135_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_136_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_137_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_138_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_139_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_140_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_141_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_142_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_143_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_144_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_145_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_146_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_147_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_148_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_149_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_150_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_151_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_152_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_153_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_154_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_155_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_156_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_157_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_158_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_159_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_160_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_161_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_162_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_163_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_164_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_165_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_166_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_167_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_168_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_169_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_170_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_171_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_172_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_173_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_174_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_175_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_176_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_177_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_178_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_179_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_180_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_181_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_182_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_183_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_184_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_185_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_186_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_187_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_188_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_189_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_190_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_191_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_192_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_193_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_194_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_195_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_196_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_197_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_198_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_199_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_200_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_201_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_202_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_203_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_204_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_205_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_206_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_207_final_cword;
