              flogtanh0xffffffff_0 = 
          (!flogtanh_sel[8]) ? 
                       flogtanh0x00008_0_q: 
                       flogtanh0x00008_1_q;
               flogtanh0xffffffff_1 =  0;
