              fgallag0x00006_0 = 
          (!fgallag_sel[5]) ? 
                       fgallag0x00005_0_q: 
                       fgallag0x00005_1_q;
              fgallag0x00006_1 = 
          (!fgallag_sel[5]) ? 
                       fgallag0x00005_2_q: 
                       fgallag0x00005_3_q;
              fgallag0x00006_2 = 
          (!fgallag_sel[5]) ? 
                       fgallag0x00005_4_q: 
                       fgallag0x00005_5_q;
              fgallag0x00006_3 = 
          (!fgallag_sel[5]) ? 
                       fgallag0x00005_6_q: 
                       fgallag0x00005_7_q;
              fgallag0x00006_4 = 
          (!fgallag_sel[5]) ? 
                       fgallag0x00005_8_q: 
                       fgallag0x00005_9_q;
              fgallag0x00006_5 = 
          (!fgallag_sel[5]) ? 
                       fgallag0x00005_10_q: 
                       fgallag0x00005_11_q;
