.o_LDPC_ENC_MSG_IN_0_msg_in(o_LDPC_ENC_MSG_IN_0_msg_in),
.o_LDPC_ENC_MSG_IN_1_msg_in(o_LDPC_ENC_MSG_IN_1_msg_in),
.o_LDPC_ENC_MSG_IN_2_msg_in(o_LDPC_ENC_MSG_IN_2_msg_in),
.o_LDPC_ENC_MSG_IN_3_msg_in(o_LDPC_ENC_MSG_IN_3_msg_in),
.o_LDPC_ENC_MSG_IN_4_msg_in(o_LDPC_ENC_MSG_IN_4_msg_in),
.o_LDPC_ENC_MSG_IN_5_msg_in(o_LDPC_ENC_MSG_IN_5_msg_in),
.o_LDPC_ENC_MSG_IN_6_msg_in(o_LDPC_ENC_MSG_IN_6_msg_in),
.o_LDPC_ENC_MSG_IN_7_msg_in(o_LDPC_ENC_MSG_IN_7_msg_in),
.o_LDPC_ENC_MSG_IN_8_msg_in(o_LDPC_ENC_MSG_IN_8_msg_in),
.o_LDPC_ENC_MSG_IN_9_msg_in(o_LDPC_ENC_MSG_IN_9_msg_in),
.o_LDPC_ENC_MSG_IN_10_msg_in(o_LDPC_ENC_MSG_IN_10_msg_in),
.o_LDPC_ENC_MSG_IN_11_msg_in(o_LDPC_ENC_MSG_IN_11_msg_in),
.o_LDPC_ENC_MSG_IN_12_msg_in(o_LDPC_ENC_MSG_IN_12_msg_in),
.o_LDPC_ENC_MSG_IN_13_msg_in(o_LDPC_ENC_MSG_IN_13_msg_in),
.o_LDPC_ENC_MSG_IN_14_msg_in(o_LDPC_ENC_MSG_IN_14_msg_in),
.o_LDPC_ENC_MSG_IN_15_msg_in(o_LDPC_ENC_MSG_IN_15_msg_in),
.o_LDPC_ENC_MSG_IN_16_msg_in(o_LDPC_ENC_MSG_IN_16_msg_in),
.o_LDPC_ENC_MSG_IN_17_msg_in(o_LDPC_ENC_MSG_IN_17_msg_in),
.o_LDPC_ENC_MSG_IN_18_msg_in(o_LDPC_ENC_MSG_IN_18_msg_in),
.o_LDPC_ENC_MSG_IN_19_msg_in(o_LDPC_ENC_MSG_IN_19_msg_in),
.o_LDPC_ENC_MSG_IN_20_msg_in(o_LDPC_ENC_MSG_IN_20_msg_in),
.o_LDPC_ENC_MSG_IN_21_msg_in(o_LDPC_ENC_MSG_IN_21_msg_in),
.o_LDPC_ENC_MSG_IN_22_msg_in(o_LDPC_ENC_MSG_IN_22_msg_in),
.o_LDPC_ENC_MSG_IN_23_msg_in(o_LDPC_ENC_MSG_IN_23_msg_in),
.o_LDPC_ENC_MSG_IN_24_msg_in(o_LDPC_ENC_MSG_IN_24_msg_in),
.o_LDPC_ENC_MSG_IN_25_msg_in(o_LDPC_ENC_MSG_IN_25_msg_in),
.o_LDPC_ENC_MSG_IN_26_msg_in(o_LDPC_ENC_MSG_IN_26_msg_in),
.o_LDPC_ENC_MSG_IN_27_msg_in(o_LDPC_ENC_MSG_IN_27_msg_in),
.o_LDPC_ENC_MSG_IN_28_msg_in(o_LDPC_ENC_MSG_IN_28_msg_in),
.o_LDPC_ENC_MSG_IN_29_msg_in(o_LDPC_ENC_MSG_IN_29_msg_in),
.o_LDPC_ENC_MSG_IN_30_msg_in(o_LDPC_ENC_MSG_IN_30_msg_in),
.o_LDPC_ENC_MSG_IN_31_msg_in(o_LDPC_ENC_MSG_IN_31_msg_in),
.o_LDPC_ENC_MSG_IN_32_msg_in(o_LDPC_ENC_MSG_IN_32_msg_in),
.o_LDPC_ENC_MSG_IN_33_msg_in(o_LDPC_ENC_MSG_IN_33_msg_in),
.o_LDPC_ENC_MSG_IN_34_msg_in(o_LDPC_ENC_MSG_IN_34_msg_in),
.o_LDPC_ENC_MSG_IN_35_msg_in(o_LDPC_ENC_MSG_IN_35_msg_in),
.o_LDPC_ENC_MSG_IN_36_msg_in(o_LDPC_ENC_MSG_IN_36_msg_in),
.o_LDPC_ENC_MSG_IN_37_msg_in(o_LDPC_ENC_MSG_IN_37_msg_in),
.o_LDPC_ENC_MSG_IN_38_msg_in(o_LDPC_ENC_MSG_IN_38_msg_in),
.o_LDPC_ENC_MSG_IN_39_msg_in(o_LDPC_ENC_MSG_IN_39_msg_in),
.i_LDPC_ENC_CODEWRD_OUT_0_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_0_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_1_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_1_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_2_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_2_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_3_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_3_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_4_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_4_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_5_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_5_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_6_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_6_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_7_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_7_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_8_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_8_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_9_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_9_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_10_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_10_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_11_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_11_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_12_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_12_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_13_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_13_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_14_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_14_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_15_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_15_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_16_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_16_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_17_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_17_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_18_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_18_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_19_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_19_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_20_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_20_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_21_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_21_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_22_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_22_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_23_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_23_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_24_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_24_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_25_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_25_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_26_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_26_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_27_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_27_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_28_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_28_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_29_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_29_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_30_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_30_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_31_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_31_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_32_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_32_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_33_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_33_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_34_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_34_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_35_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_35_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_36_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_36_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_37_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_37_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_38_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_38_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_39_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_39_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_40_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_40_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_41_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_41_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_42_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_42_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_43_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_43_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_44_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_44_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_45_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_45_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_46_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_46_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_47_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_47_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_48_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_48_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_49_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_49_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_50_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_50_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_51_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_51_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_52_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_52_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_53_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_53_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_54_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_54_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_55_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_55_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_56_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_56_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_57_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_57_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_58_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_58_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_59_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_59_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_60_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_60_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_61_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_61_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_62_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_62_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_63_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_63_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_64_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_64_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_65_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_65_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_66_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_66_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_67_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_67_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_68_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_68_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_69_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_69_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_70_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_70_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_71_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_71_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_72_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_72_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_73_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_73_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_74_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_74_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_75_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_75_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_76_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_76_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_77_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_77_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_78_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_78_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_79_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_79_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_80_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_80_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_81_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_81_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_82_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_82_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_83_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_83_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_84_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_84_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_85_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_85_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_86_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_86_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_87_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_87_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_88_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_88_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_89_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_89_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_90_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_90_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_91_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_91_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_92_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_92_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_93_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_93_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_94_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_94_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_95_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_95_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_96_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_96_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_97_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_97_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_98_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_98_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_99_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_99_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_100_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_100_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_101_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_101_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_102_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_102_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_103_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_103_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_104_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_104_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_105_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_105_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_106_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_106_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_107_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_107_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_108_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_108_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_109_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_109_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_110_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_110_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_111_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_111_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_112_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_112_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_113_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_113_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_114_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_114_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_115_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_115_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_116_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_116_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_117_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_117_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_118_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_118_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_119_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_119_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_120_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_120_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_121_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_121_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_122_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_122_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_123_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_123_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_124_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_124_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_125_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_125_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_126_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_126_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_127_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_127_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_128_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_128_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_129_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_129_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_130_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_130_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_131_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_131_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_132_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_132_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_133_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_133_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_134_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_134_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_135_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_135_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_136_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_136_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_137_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_137_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_138_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_138_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_139_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_139_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_140_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_140_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_141_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_141_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_142_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_142_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_143_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_143_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_144_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_144_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_145_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_145_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_146_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_146_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_147_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_147_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_148_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_148_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_149_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_149_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_150_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_150_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_151_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_151_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_152_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_152_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_153_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_153_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_154_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_154_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_155_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_155_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_156_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_156_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_157_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_157_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_158_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_158_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_159_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_159_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_160_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_160_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_161_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_161_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_162_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_162_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_163_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_163_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_164_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_164_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_165_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_165_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_166_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_166_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_167_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_167_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_168_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_168_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_169_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_169_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_170_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_170_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_171_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_171_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_172_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_172_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_173_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_173_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_174_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_174_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_175_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_175_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_176_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_176_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_177_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_177_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_178_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_178_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_179_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_179_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_180_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_180_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_181_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_181_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_182_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_182_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_183_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_183_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_184_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_184_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_185_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_185_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_186_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_186_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_187_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_187_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_188_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_188_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_189_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_189_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_190_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_190_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_191_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_191_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_192_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_192_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_193_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_193_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_194_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_194_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_195_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_195_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_196_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_196_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_197_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_197_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_198_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_198_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_199_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_199_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_200_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_200_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_201_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_201_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_202_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_202_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_203_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_203_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_204_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_204_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_205_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_205_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_206_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_206_enc_codeword),
.i_LDPC_ENC_CODEWRD_OUT_207_enc_codeword(i_LDPC_ENC_CODEWRD_OUT_207_enc_codeword),
.i_LDPC_ENC_CODEWRD_VLD_enc_codeword_valid(i_LDPC_ENC_CODEWRD_VLD_enc_codeword_valid),
.o_LDPC_DEC_ERR_INTRODUCED_err_intro(o_LDPC_DEC_ERR_INTRODUCED_err_intro),
.o_LDPC_DEC_SEL_FRMC_sel_q0_frmC(o_LDPC_DEC_SEL_FRMC_sel_q0_frmC),
.o_LDPC_DEC_ERR_Q0_0_INTRO_0_err_intro_q0_0_0(o_LDPC_DEC_ERR_Q0_0_INTRO_0_err_intro_q0_0_0),
.o_LDPC_DEC_ERR_Q0_0_INTRO_1_err_intro_q0_0_1(o_LDPC_DEC_ERR_Q0_0_INTRO_1_err_intro_q0_0_1),
.o_LDPC_DEC_ERR_Q0_0_INTRO_2_err_intro_q0_0_2(o_LDPC_DEC_ERR_Q0_0_INTRO_2_err_intro_q0_0_2),
.o_LDPC_DEC_ERR_Q0_0_INTRO_3_err_intro_q0_0_3(o_LDPC_DEC_ERR_Q0_0_INTRO_3_err_intro_q0_0_3),
.o_LDPC_DEC_ERR_Q0_0_INTRO_4_err_intro_q0_0_4(o_LDPC_DEC_ERR_Q0_0_INTRO_4_err_intro_q0_0_4),
.o_LDPC_DEC_ERR_Q0_0_INTRO_5_err_intro_q0_0_5(o_LDPC_DEC_ERR_Q0_0_INTRO_5_err_intro_q0_0_5),
.o_LDPC_DEC_ERR_Q0_0_INTRO_6_err_intro_q0_0_6(o_LDPC_DEC_ERR_Q0_0_INTRO_6_err_intro_q0_0_6),
.o_LDPC_DEC_ERR_Q0_0_INTRO_7_err_intro_q0_0_7(o_LDPC_DEC_ERR_Q0_0_INTRO_7_err_intro_q0_0_7),
.o_LDPC_DEC_ERR_Q0_0_INTRO_8_err_intro_q0_0_8(o_LDPC_DEC_ERR_Q0_0_INTRO_8_err_intro_q0_0_8),
.o_LDPC_DEC_ERR_Q0_0_INTRO_9_err_intro_q0_0_9(o_LDPC_DEC_ERR_Q0_0_INTRO_9_err_intro_q0_0_9),
.o_LDPC_DEC_ERR_Q0_0_INTRO_10_err_intro_q0_0_10(o_LDPC_DEC_ERR_Q0_0_INTRO_10_err_intro_q0_0_10),
.o_LDPC_DEC_ERR_Q0_0_INTRO_11_err_intro_q0_0_11(o_LDPC_DEC_ERR_Q0_0_INTRO_11_err_intro_q0_0_11),
.o_LDPC_DEC_ERR_Q0_0_INTRO_12_err_intro_q0_0_12(o_LDPC_DEC_ERR_Q0_0_INTRO_12_err_intro_q0_0_12),
.o_LDPC_DEC_ERR_Q0_0_INTRO_13_err_intro_q0_0_13(o_LDPC_DEC_ERR_Q0_0_INTRO_13_err_intro_q0_0_13),
.o_LDPC_DEC_ERR_Q0_0_INTRO_14_err_intro_q0_0_14(o_LDPC_DEC_ERR_Q0_0_INTRO_14_err_intro_q0_0_14),
.o_LDPC_DEC_ERR_Q0_0_INTRO_15_err_intro_q0_0_15(o_LDPC_DEC_ERR_Q0_0_INTRO_15_err_intro_q0_0_15),
.o_LDPC_DEC_ERR_Q0_0_INTRO_16_err_intro_q0_0_16(o_LDPC_DEC_ERR_Q0_0_INTRO_16_err_intro_q0_0_16),
.o_LDPC_DEC_ERR_Q0_0_INTRO_17_err_intro_q0_0_17(o_LDPC_DEC_ERR_Q0_0_INTRO_17_err_intro_q0_0_17),
.o_LDPC_DEC_ERR_Q0_0_INTRO_18_err_intro_q0_0_18(o_LDPC_DEC_ERR_Q0_0_INTRO_18_err_intro_q0_0_18),
.o_LDPC_DEC_ERR_Q0_0_INTRO_19_err_intro_q0_0_19(o_LDPC_DEC_ERR_Q0_0_INTRO_19_err_intro_q0_0_19),
.o_LDPC_DEC_ERR_Q0_0_INTRO_20_err_intro_q0_0_20(o_LDPC_DEC_ERR_Q0_0_INTRO_20_err_intro_q0_0_20),
.o_LDPC_DEC_ERR_Q0_0_INTRO_21_err_intro_q0_0_21(o_LDPC_DEC_ERR_Q0_0_INTRO_21_err_intro_q0_0_21),
.o_LDPC_DEC_ERR_Q0_0_INTRO_22_err_intro_q0_0_22(o_LDPC_DEC_ERR_Q0_0_INTRO_22_err_intro_q0_0_22),
.o_LDPC_DEC_ERR_Q0_0_INTRO_23_err_intro_q0_0_23(o_LDPC_DEC_ERR_Q0_0_INTRO_23_err_intro_q0_0_23),
.o_LDPC_DEC_ERR_Q0_0_INTRO_24_err_intro_q0_0_24(o_LDPC_DEC_ERR_Q0_0_INTRO_24_err_intro_q0_0_24),
.o_LDPC_DEC_ERR_Q0_0_INTRO_25_err_intro_q0_0_25(o_LDPC_DEC_ERR_Q0_0_INTRO_25_err_intro_q0_0_25),
.o_LDPC_DEC_ERR_Q0_0_INTRO_26_err_intro_q0_0_26(o_LDPC_DEC_ERR_Q0_0_INTRO_26_err_intro_q0_0_26),
.o_LDPC_DEC_ERR_Q0_0_INTRO_27_err_intro_q0_0_27(o_LDPC_DEC_ERR_Q0_0_INTRO_27_err_intro_q0_0_27),
.o_LDPC_DEC_ERR_Q0_0_INTRO_28_err_intro_q0_0_28(o_LDPC_DEC_ERR_Q0_0_INTRO_28_err_intro_q0_0_28),
.o_LDPC_DEC_ERR_Q0_0_INTRO_29_err_intro_q0_0_29(o_LDPC_DEC_ERR_Q0_0_INTRO_29_err_intro_q0_0_29),
.o_LDPC_DEC_ERR_Q0_0_INTRO_30_err_intro_q0_0_30(o_LDPC_DEC_ERR_Q0_0_INTRO_30_err_intro_q0_0_30),
.o_LDPC_DEC_ERR_Q0_0_INTRO_31_err_intro_q0_0_31(o_LDPC_DEC_ERR_Q0_0_INTRO_31_err_intro_q0_0_31),
.o_LDPC_DEC_ERR_Q0_0_INTRO_32_err_intro_q0_0_32(o_LDPC_DEC_ERR_Q0_0_INTRO_32_err_intro_q0_0_32),
.o_LDPC_DEC_ERR_Q0_0_INTRO_33_err_intro_q0_0_33(o_LDPC_DEC_ERR_Q0_0_INTRO_33_err_intro_q0_0_33),
.o_LDPC_DEC_ERR_Q0_0_INTRO_34_err_intro_q0_0_34(o_LDPC_DEC_ERR_Q0_0_INTRO_34_err_intro_q0_0_34),
.o_LDPC_DEC_ERR_Q0_0_INTRO_35_err_intro_q0_0_35(o_LDPC_DEC_ERR_Q0_0_INTRO_35_err_intro_q0_0_35),
.o_LDPC_DEC_ERR_Q0_0_INTRO_36_err_intro_q0_0_36(o_LDPC_DEC_ERR_Q0_0_INTRO_36_err_intro_q0_0_36),
.o_LDPC_DEC_ERR_Q0_0_INTRO_37_err_intro_q0_0_37(o_LDPC_DEC_ERR_Q0_0_INTRO_37_err_intro_q0_0_37),
.o_LDPC_DEC_ERR_Q0_0_INTRO_38_err_intro_q0_0_38(o_LDPC_DEC_ERR_Q0_0_INTRO_38_err_intro_q0_0_38),
.o_LDPC_DEC_ERR_Q0_0_INTRO_39_err_intro_q0_0_39(o_LDPC_DEC_ERR_Q0_0_INTRO_39_err_intro_q0_0_39),
.o_LDPC_DEC_ERR_Q0_0_INTRO_40_err_intro_q0_0_40(o_LDPC_DEC_ERR_Q0_0_INTRO_40_err_intro_q0_0_40),
.o_LDPC_DEC_ERR_Q0_0_INTRO_41_err_intro_q0_0_41(o_LDPC_DEC_ERR_Q0_0_INTRO_41_err_intro_q0_0_41),
.o_LDPC_DEC_ERR_Q0_0_INTRO_42_err_intro_q0_0_42(o_LDPC_DEC_ERR_Q0_0_INTRO_42_err_intro_q0_0_42),
.o_LDPC_DEC_ERR_Q0_0_INTRO_43_err_intro_q0_0_43(o_LDPC_DEC_ERR_Q0_0_INTRO_43_err_intro_q0_0_43),
.o_LDPC_DEC_ERR_Q0_0_INTRO_44_err_intro_q0_0_44(o_LDPC_DEC_ERR_Q0_0_INTRO_44_err_intro_q0_0_44),
.o_LDPC_DEC_ERR_Q0_0_INTRO_45_err_intro_q0_0_45(o_LDPC_DEC_ERR_Q0_0_INTRO_45_err_intro_q0_0_45),
.o_LDPC_DEC_ERR_Q0_0_INTRO_46_err_intro_q0_0_46(o_LDPC_DEC_ERR_Q0_0_INTRO_46_err_intro_q0_0_46),
.o_LDPC_DEC_ERR_Q0_0_INTRO_47_err_intro_q0_0_47(o_LDPC_DEC_ERR_Q0_0_INTRO_47_err_intro_q0_0_47),
.o_LDPC_DEC_ERR_Q0_0_INTRO_48_err_intro_q0_0_48(o_LDPC_DEC_ERR_Q0_0_INTRO_48_err_intro_q0_0_48),
.o_LDPC_DEC_ERR_Q0_0_INTRO_49_err_intro_q0_0_49(o_LDPC_DEC_ERR_Q0_0_INTRO_49_err_intro_q0_0_49),
.o_LDPC_DEC_ERR_Q0_0_INTRO_50_err_intro_q0_0_50(o_LDPC_DEC_ERR_Q0_0_INTRO_50_err_intro_q0_0_50),
.o_LDPC_DEC_ERR_Q0_0_INTRO_51_err_intro_q0_0_51(o_LDPC_DEC_ERR_Q0_0_INTRO_51_err_intro_q0_0_51),
.o_LDPC_DEC_ERR_Q0_0_INTRO_52_err_intro_q0_0_52(o_LDPC_DEC_ERR_Q0_0_INTRO_52_err_intro_q0_0_52),
.o_LDPC_DEC_ERR_Q0_0_INTRO_53_err_intro_q0_0_53(o_LDPC_DEC_ERR_Q0_0_INTRO_53_err_intro_q0_0_53),
.o_LDPC_DEC_ERR_Q0_0_INTRO_54_err_intro_q0_0_54(o_LDPC_DEC_ERR_Q0_0_INTRO_54_err_intro_q0_0_54),
.o_LDPC_DEC_ERR_Q0_0_INTRO_55_err_intro_q0_0_55(o_LDPC_DEC_ERR_Q0_0_INTRO_55_err_intro_q0_0_55),
.o_LDPC_DEC_ERR_Q0_0_INTRO_56_err_intro_q0_0_56(o_LDPC_DEC_ERR_Q0_0_INTRO_56_err_intro_q0_0_56),
.o_LDPC_DEC_ERR_Q0_0_INTRO_57_err_intro_q0_0_57(o_LDPC_DEC_ERR_Q0_0_INTRO_57_err_intro_q0_0_57),
.o_LDPC_DEC_ERR_Q0_0_INTRO_58_err_intro_q0_0_58(o_LDPC_DEC_ERR_Q0_0_INTRO_58_err_intro_q0_0_58),
.o_LDPC_DEC_ERR_Q0_0_INTRO_59_err_intro_q0_0_59(o_LDPC_DEC_ERR_Q0_0_INTRO_59_err_intro_q0_0_59),
.o_LDPC_DEC_ERR_Q0_0_INTRO_60_err_intro_q0_0_60(o_LDPC_DEC_ERR_Q0_0_INTRO_60_err_intro_q0_0_60),
.o_LDPC_DEC_ERR_Q0_0_INTRO_61_err_intro_q0_0_61(o_LDPC_DEC_ERR_Q0_0_INTRO_61_err_intro_q0_0_61),
.o_LDPC_DEC_ERR_Q0_0_INTRO_62_err_intro_q0_0_62(o_LDPC_DEC_ERR_Q0_0_INTRO_62_err_intro_q0_0_62),
.o_LDPC_DEC_ERR_Q0_0_INTRO_63_err_intro_q0_0_63(o_LDPC_DEC_ERR_Q0_0_INTRO_63_err_intro_q0_0_63),
.o_LDPC_DEC_ERR_Q0_0_INTRO_64_err_intro_q0_0_64(o_LDPC_DEC_ERR_Q0_0_INTRO_64_err_intro_q0_0_64),
.o_LDPC_DEC_ERR_Q0_0_INTRO_65_err_intro_q0_0_65(o_LDPC_DEC_ERR_Q0_0_INTRO_65_err_intro_q0_0_65),
.o_LDPC_DEC_ERR_Q0_0_INTRO_66_err_intro_q0_0_66(o_LDPC_DEC_ERR_Q0_0_INTRO_66_err_intro_q0_0_66),
.o_LDPC_DEC_ERR_Q0_0_INTRO_67_err_intro_q0_0_67(o_LDPC_DEC_ERR_Q0_0_INTRO_67_err_intro_q0_0_67),
.o_LDPC_DEC_ERR_Q0_0_INTRO_68_err_intro_q0_0_68(o_LDPC_DEC_ERR_Q0_0_INTRO_68_err_intro_q0_0_68),
.o_LDPC_DEC_ERR_Q0_0_INTRO_69_err_intro_q0_0_69(o_LDPC_DEC_ERR_Q0_0_INTRO_69_err_intro_q0_0_69),
.o_LDPC_DEC_ERR_Q0_0_INTRO_70_err_intro_q0_0_70(o_LDPC_DEC_ERR_Q0_0_INTRO_70_err_intro_q0_0_70),
.o_LDPC_DEC_ERR_Q0_0_INTRO_71_err_intro_q0_0_71(o_LDPC_DEC_ERR_Q0_0_INTRO_71_err_intro_q0_0_71),
.o_LDPC_DEC_ERR_Q0_0_INTRO_72_err_intro_q0_0_72(o_LDPC_DEC_ERR_Q0_0_INTRO_72_err_intro_q0_0_72),
.o_LDPC_DEC_ERR_Q0_0_INTRO_73_err_intro_q0_0_73(o_LDPC_DEC_ERR_Q0_0_INTRO_73_err_intro_q0_0_73),
.o_LDPC_DEC_ERR_Q0_0_INTRO_74_err_intro_q0_0_74(o_LDPC_DEC_ERR_Q0_0_INTRO_74_err_intro_q0_0_74),
.o_LDPC_DEC_ERR_Q0_0_INTRO_75_err_intro_q0_0_75(o_LDPC_DEC_ERR_Q0_0_INTRO_75_err_intro_q0_0_75),
.o_LDPC_DEC_ERR_Q0_0_INTRO_76_err_intro_q0_0_76(o_LDPC_DEC_ERR_Q0_0_INTRO_76_err_intro_q0_0_76),
.o_LDPC_DEC_ERR_Q0_0_INTRO_77_err_intro_q0_0_77(o_LDPC_DEC_ERR_Q0_0_INTRO_77_err_intro_q0_0_77),
.o_LDPC_DEC_ERR_Q0_0_INTRO_78_err_intro_q0_0_78(o_LDPC_DEC_ERR_Q0_0_INTRO_78_err_intro_q0_0_78),
.o_LDPC_DEC_ERR_Q0_0_INTRO_79_err_intro_q0_0_79(o_LDPC_DEC_ERR_Q0_0_INTRO_79_err_intro_q0_0_79),
.o_LDPC_DEC_ERR_Q0_0_INTRO_80_err_intro_q0_0_80(o_LDPC_DEC_ERR_Q0_0_INTRO_80_err_intro_q0_0_80),
.o_LDPC_DEC_ERR_Q0_0_INTRO_81_err_intro_q0_0_81(o_LDPC_DEC_ERR_Q0_0_INTRO_81_err_intro_q0_0_81),
.o_LDPC_DEC_ERR_Q0_0_INTRO_82_err_intro_q0_0_82(o_LDPC_DEC_ERR_Q0_0_INTRO_82_err_intro_q0_0_82),
.o_LDPC_DEC_ERR_Q0_0_INTRO_83_err_intro_q0_0_83(o_LDPC_DEC_ERR_Q0_0_INTRO_83_err_intro_q0_0_83),
.o_LDPC_DEC_ERR_Q0_0_INTRO_84_err_intro_q0_0_84(o_LDPC_DEC_ERR_Q0_0_INTRO_84_err_intro_q0_0_84),
.o_LDPC_DEC_ERR_Q0_0_INTRO_85_err_intro_q0_0_85(o_LDPC_DEC_ERR_Q0_0_INTRO_85_err_intro_q0_0_85),
.o_LDPC_DEC_ERR_Q0_0_INTRO_86_err_intro_q0_0_86(o_LDPC_DEC_ERR_Q0_0_INTRO_86_err_intro_q0_0_86),
.o_LDPC_DEC_ERR_Q0_0_INTRO_87_err_intro_q0_0_87(o_LDPC_DEC_ERR_Q0_0_INTRO_87_err_intro_q0_0_87),
.o_LDPC_DEC_ERR_Q0_0_INTRO_88_err_intro_q0_0_88(o_LDPC_DEC_ERR_Q0_0_INTRO_88_err_intro_q0_0_88),
.o_LDPC_DEC_ERR_Q0_0_INTRO_89_err_intro_q0_0_89(o_LDPC_DEC_ERR_Q0_0_INTRO_89_err_intro_q0_0_89),
.o_LDPC_DEC_ERR_Q0_0_INTRO_90_err_intro_q0_0_90(o_LDPC_DEC_ERR_Q0_0_INTRO_90_err_intro_q0_0_90),
.o_LDPC_DEC_ERR_Q0_0_INTRO_91_err_intro_q0_0_91(o_LDPC_DEC_ERR_Q0_0_INTRO_91_err_intro_q0_0_91),
.o_LDPC_DEC_ERR_Q0_0_INTRO_92_err_intro_q0_0_92(o_LDPC_DEC_ERR_Q0_0_INTRO_92_err_intro_q0_0_92),
.o_LDPC_DEC_ERR_Q0_0_INTRO_93_err_intro_q0_0_93(o_LDPC_DEC_ERR_Q0_0_INTRO_93_err_intro_q0_0_93),
.o_LDPC_DEC_ERR_Q0_0_INTRO_94_err_intro_q0_0_94(o_LDPC_DEC_ERR_Q0_0_INTRO_94_err_intro_q0_0_94),
.o_LDPC_DEC_ERR_Q0_0_INTRO_95_err_intro_q0_0_95(o_LDPC_DEC_ERR_Q0_0_INTRO_95_err_intro_q0_0_95),
.o_LDPC_DEC_ERR_Q0_0_INTRO_96_err_intro_q0_0_96(o_LDPC_DEC_ERR_Q0_0_INTRO_96_err_intro_q0_0_96),
.o_LDPC_DEC_ERR_Q0_0_INTRO_97_err_intro_q0_0_97(o_LDPC_DEC_ERR_Q0_0_INTRO_97_err_intro_q0_0_97),
.o_LDPC_DEC_ERR_Q0_0_INTRO_98_err_intro_q0_0_98(o_LDPC_DEC_ERR_Q0_0_INTRO_98_err_intro_q0_0_98),
.o_LDPC_DEC_ERR_Q0_0_INTRO_99_err_intro_q0_0_99(o_LDPC_DEC_ERR_Q0_0_INTRO_99_err_intro_q0_0_99),
.o_LDPC_DEC_ERR_Q0_0_INTRO_100_err_intro_q0_0_100(o_LDPC_DEC_ERR_Q0_0_INTRO_100_err_intro_q0_0_100),
.o_LDPC_DEC_ERR_Q0_0_INTRO_101_err_intro_q0_0_101(o_LDPC_DEC_ERR_Q0_0_INTRO_101_err_intro_q0_0_101),
.o_LDPC_DEC_ERR_Q0_0_INTRO_102_err_intro_q0_0_102(o_LDPC_DEC_ERR_Q0_0_INTRO_102_err_intro_q0_0_102),
.o_LDPC_DEC_ERR_Q0_0_INTRO_103_err_intro_q0_0_103(o_LDPC_DEC_ERR_Q0_0_INTRO_103_err_intro_q0_0_103),
.o_LDPC_DEC_ERR_Q0_0_INTRO_104_err_intro_q0_0_104(o_LDPC_DEC_ERR_Q0_0_INTRO_104_err_intro_q0_0_104),
.o_LDPC_DEC_ERR_Q0_0_INTRO_105_err_intro_q0_0_105(o_LDPC_DEC_ERR_Q0_0_INTRO_105_err_intro_q0_0_105),
.o_LDPC_DEC_ERR_Q0_0_INTRO_106_err_intro_q0_0_106(o_LDPC_DEC_ERR_Q0_0_INTRO_106_err_intro_q0_0_106),
.o_LDPC_DEC_ERR_Q0_0_INTRO_107_err_intro_q0_0_107(o_LDPC_DEC_ERR_Q0_0_INTRO_107_err_intro_q0_0_107),
.o_LDPC_DEC_ERR_Q0_0_INTRO_108_err_intro_q0_0_108(o_LDPC_DEC_ERR_Q0_0_INTRO_108_err_intro_q0_0_108),
.o_LDPC_DEC_ERR_Q0_0_INTRO_109_err_intro_q0_0_109(o_LDPC_DEC_ERR_Q0_0_INTRO_109_err_intro_q0_0_109),
.o_LDPC_DEC_ERR_Q0_0_INTRO_110_err_intro_q0_0_110(o_LDPC_DEC_ERR_Q0_0_INTRO_110_err_intro_q0_0_110),
.o_LDPC_DEC_ERR_Q0_0_INTRO_111_err_intro_q0_0_111(o_LDPC_DEC_ERR_Q0_0_INTRO_111_err_intro_q0_0_111),
.o_LDPC_DEC_ERR_Q0_0_INTRO_112_err_intro_q0_0_112(o_LDPC_DEC_ERR_Q0_0_INTRO_112_err_intro_q0_0_112),
.o_LDPC_DEC_ERR_Q0_0_INTRO_113_err_intro_q0_0_113(o_LDPC_DEC_ERR_Q0_0_INTRO_113_err_intro_q0_0_113),
.o_LDPC_DEC_ERR_Q0_0_INTRO_114_err_intro_q0_0_114(o_LDPC_DEC_ERR_Q0_0_INTRO_114_err_intro_q0_0_114),
.o_LDPC_DEC_ERR_Q0_0_INTRO_115_err_intro_q0_0_115(o_LDPC_DEC_ERR_Q0_0_INTRO_115_err_intro_q0_0_115),
.o_LDPC_DEC_ERR_Q0_0_INTRO_116_err_intro_q0_0_116(o_LDPC_DEC_ERR_Q0_0_INTRO_116_err_intro_q0_0_116),
.o_LDPC_DEC_ERR_Q0_0_INTRO_117_err_intro_q0_0_117(o_LDPC_DEC_ERR_Q0_0_INTRO_117_err_intro_q0_0_117),
.o_LDPC_DEC_ERR_Q0_0_INTRO_118_err_intro_q0_0_118(o_LDPC_DEC_ERR_Q0_0_INTRO_118_err_intro_q0_0_118),
.o_LDPC_DEC_ERR_Q0_0_INTRO_119_err_intro_q0_0_119(o_LDPC_DEC_ERR_Q0_0_INTRO_119_err_intro_q0_0_119),
.o_LDPC_DEC_ERR_Q0_0_INTRO_120_err_intro_q0_0_120(o_LDPC_DEC_ERR_Q0_0_INTRO_120_err_intro_q0_0_120),
.o_LDPC_DEC_ERR_Q0_0_INTRO_121_err_intro_q0_0_121(o_LDPC_DEC_ERR_Q0_0_INTRO_121_err_intro_q0_0_121),
.o_LDPC_DEC_ERR_Q0_0_INTRO_122_err_intro_q0_0_122(o_LDPC_DEC_ERR_Q0_0_INTRO_122_err_intro_q0_0_122),
.o_LDPC_DEC_ERR_Q0_0_INTRO_123_err_intro_q0_0_123(o_LDPC_DEC_ERR_Q0_0_INTRO_123_err_intro_q0_0_123),
.o_LDPC_DEC_ERR_Q0_0_INTRO_124_err_intro_q0_0_124(o_LDPC_DEC_ERR_Q0_0_INTRO_124_err_intro_q0_0_124),
.o_LDPC_DEC_ERR_Q0_0_INTRO_125_err_intro_q0_0_125(o_LDPC_DEC_ERR_Q0_0_INTRO_125_err_intro_q0_0_125),
.o_LDPC_DEC_ERR_Q0_0_INTRO_126_err_intro_q0_0_126(o_LDPC_DEC_ERR_Q0_0_INTRO_126_err_intro_q0_0_126),
.o_LDPC_DEC_ERR_Q0_0_INTRO_127_err_intro_q0_0_127(o_LDPC_DEC_ERR_Q0_0_INTRO_127_err_intro_q0_0_127),
.o_LDPC_DEC_ERR_Q0_0_INTRO_128_err_intro_q0_0_128(o_LDPC_DEC_ERR_Q0_0_INTRO_128_err_intro_q0_0_128),
.o_LDPC_DEC_ERR_Q0_0_INTRO_129_err_intro_q0_0_129(o_LDPC_DEC_ERR_Q0_0_INTRO_129_err_intro_q0_0_129),
.o_LDPC_DEC_ERR_Q0_0_INTRO_130_err_intro_q0_0_130(o_LDPC_DEC_ERR_Q0_0_INTRO_130_err_intro_q0_0_130),
.o_LDPC_DEC_ERR_Q0_0_INTRO_131_err_intro_q0_0_131(o_LDPC_DEC_ERR_Q0_0_INTRO_131_err_intro_q0_0_131),
.o_LDPC_DEC_ERR_Q0_0_INTRO_132_err_intro_q0_0_132(o_LDPC_DEC_ERR_Q0_0_INTRO_132_err_intro_q0_0_132),
.o_LDPC_DEC_ERR_Q0_0_INTRO_133_err_intro_q0_0_133(o_LDPC_DEC_ERR_Q0_0_INTRO_133_err_intro_q0_0_133),
.o_LDPC_DEC_ERR_Q0_0_INTRO_134_err_intro_q0_0_134(o_LDPC_DEC_ERR_Q0_0_INTRO_134_err_intro_q0_0_134),
.o_LDPC_DEC_ERR_Q0_0_INTRO_135_err_intro_q0_0_135(o_LDPC_DEC_ERR_Q0_0_INTRO_135_err_intro_q0_0_135),
.o_LDPC_DEC_ERR_Q0_0_INTRO_136_err_intro_q0_0_136(o_LDPC_DEC_ERR_Q0_0_INTRO_136_err_intro_q0_0_136),
.o_LDPC_DEC_ERR_Q0_0_INTRO_137_err_intro_q0_0_137(o_LDPC_DEC_ERR_Q0_0_INTRO_137_err_intro_q0_0_137),
.o_LDPC_DEC_ERR_Q0_0_INTRO_138_err_intro_q0_0_138(o_LDPC_DEC_ERR_Q0_0_INTRO_138_err_intro_q0_0_138),
.o_LDPC_DEC_ERR_Q0_0_INTRO_139_err_intro_q0_0_139(o_LDPC_DEC_ERR_Q0_0_INTRO_139_err_intro_q0_0_139),
.o_LDPC_DEC_ERR_Q0_0_INTRO_140_err_intro_q0_0_140(o_LDPC_DEC_ERR_Q0_0_INTRO_140_err_intro_q0_0_140),
.o_LDPC_DEC_ERR_Q0_0_INTRO_141_err_intro_q0_0_141(o_LDPC_DEC_ERR_Q0_0_INTRO_141_err_intro_q0_0_141),
.o_LDPC_DEC_ERR_Q0_0_INTRO_142_err_intro_q0_0_142(o_LDPC_DEC_ERR_Q0_0_INTRO_142_err_intro_q0_0_142),
.o_LDPC_DEC_ERR_Q0_0_INTRO_143_err_intro_q0_0_143(o_LDPC_DEC_ERR_Q0_0_INTRO_143_err_intro_q0_0_143),
.o_LDPC_DEC_ERR_Q0_0_INTRO_144_err_intro_q0_0_144(o_LDPC_DEC_ERR_Q0_0_INTRO_144_err_intro_q0_0_144),
.o_LDPC_DEC_ERR_Q0_0_INTRO_145_err_intro_q0_0_145(o_LDPC_DEC_ERR_Q0_0_INTRO_145_err_intro_q0_0_145),
.o_LDPC_DEC_ERR_Q0_0_INTRO_146_err_intro_q0_0_146(o_LDPC_DEC_ERR_Q0_0_INTRO_146_err_intro_q0_0_146),
.o_LDPC_DEC_ERR_Q0_0_INTRO_147_err_intro_q0_0_147(o_LDPC_DEC_ERR_Q0_0_INTRO_147_err_intro_q0_0_147),
.o_LDPC_DEC_ERR_Q0_0_INTRO_148_err_intro_q0_0_148(o_LDPC_DEC_ERR_Q0_0_INTRO_148_err_intro_q0_0_148),
.o_LDPC_DEC_ERR_Q0_0_INTRO_149_err_intro_q0_0_149(o_LDPC_DEC_ERR_Q0_0_INTRO_149_err_intro_q0_0_149),
.o_LDPC_DEC_ERR_Q0_0_INTRO_150_err_intro_q0_0_150(o_LDPC_DEC_ERR_Q0_0_INTRO_150_err_intro_q0_0_150),
.o_LDPC_DEC_ERR_Q0_0_INTRO_151_err_intro_q0_0_151(o_LDPC_DEC_ERR_Q0_0_INTRO_151_err_intro_q0_0_151),
.o_LDPC_DEC_ERR_Q0_0_INTRO_152_err_intro_q0_0_152(o_LDPC_DEC_ERR_Q0_0_INTRO_152_err_intro_q0_0_152),
.o_LDPC_DEC_ERR_Q0_0_INTRO_153_err_intro_q0_0_153(o_LDPC_DEC_ERR_Q0_0_INTRO_153_err_intro_q0_0_153),
.o_LDPC_DEC_ERR_Q0_0_INTRO_154_err_intro_q0_0_154(o_LDPC_DEC_ERR_Q0_0_INTRO_154_err_intro_q0_0_154),
.o_LDPC_DEC_ERR_Q0_0_INTRO_155_err_intro_q0_0_155(o_LDPC_DEC_ERR_Q0_0_INTRO_155_err_intro_q0_0_155),
.o_LDPC_DEC_ERR_Q0_0_INTRO_156_err_intro_q0_0_156(o_LDPC_DEC_ERR_Q0_0_INTRO_156_err_intro_q0_0_156),
.o_LDPC_DEC_ERR_Q0_0_INTRO_157_err_intro_q0_0_157(o_LDPC_DEC_ERR_Q0_0_INTRO_157_err_intro_q0_0_157),
.o_LDPC_DEC_ERR_Q0_0_INTRO_158_err_intro_q0_0_158(o_LDPC_DEC_ERR_Q0_0_INTRO_158_err_intro_q0_0_158),
.o_LDPC_DEC_ERR_Q0_0_INTRO_159_err_intro_q0_0_159(o_LDPC_DEC_ERR_Q0_0_INTRO_159_err_intro_q0_0_159),
.o_LDPC_DEC_ERR_Q0_0_INTRO_160_err_intro_q0_0_160(o_LDPC_DEC_ERR_Q0_0_INTRO_160_err_intro_q0_0_160),
.o_LDPC_DEC_ERR_Q0_0_INTRO_161_err_intro_q0_0_161(o_LDPC_DEC_ERR_Q0_0_INTRO_161_err_intro_q0_0_161),
.o_LDPC_DEC_ERR_Q0_0_INTRO_162_err_intro_q0_0_162(o_LDPC_DEC_ERR_Q0_0_INTRO_162_err_intro_q0_0_162),
.o_LDPC_DEC_ERR_Q0_0_INTRO_163_err_intro_q0_0_163(o_LDPC_DEC_ERR_Q0_0_INTRO_163_err_intro_q0_0_163),
.o_LDPC_DEC_ERR_Q0_0_INTRO_164_err_intro_q0_0_164(o_LDPC_DEC_ERR_Q0_0_INTRO_164_err_intro_q0_0_164),
.o_LDPC_DEC_ERR_Q0_0_INTRO_165_err_intro_q0_0_165(o_LDPC_DEC_ERR_Q0_0_INTRO_165_err_intro_q0_0_165),
.o_LDPC_DEC_ERR_Q0_0_INTRO_166_err_intro_q0_0_166(o_LDPC_DEC_ERR_Q0_0_INTRO_166_err_intro_q0_0_166),
.o_LDPC_DEC_ERR_Q0_0_INTRO_167_err_intro_q0_0_167(o_LDPC_DEC_ERR_Q0_0_INTRO_167_err_intro_q0_0_167),
.o_LDPC_DEC_ERR_Q0_0_INTRO_168_err_intro_q0_0_168(o_LDPC_DEC_ERR_Q0_0_INTRO_168_err_intro_q0_0_168),
.o_LDPC_DEC_ERR_Q0_0_INTRO_169_err_intro_q0_0_169(o_LDPC_DEC_ERR_Q0_0_INTRO_169_err_intro_q0_0_169),
.o_LDPC_DEC_ERR_Q0_0_INTRO_170_err_intro_q0_0_170(o_LDPC_DEC_ERR_Q0_0_INTRO_170_err_intro_q0_0_170),
.o_LDPC_DEC_ERR_Q0_0_INTRO_171_err_intro_q0_0_171(o_LDPC_DEC_ERR_Q0_0_INTRO_171_err_intro_q0_0_171),
.o_LDPC_DEC_ERR_Q0_0_INTRO_172_err_intro_q0_0_172(o_LDPC_DEC_ERR_Q0_0_INTRO_172_err_intro_q0_0_172),
.o_LDPC_DEC_ERR_Q0_0_INTRO_173_err_intro_q0_0_173(o_LDPC_DEC_ERR_Q0_0_INTRO_173_err_intro_q0_0_173),
.o_LDPC_DEC_ERR_Q0_0_INTRO_174_err_intro_q0_0_174(o_LDPC_DEC_ERR_Q0_0_INTRO_174_err_intro_q0_0_174),
.o_LDPC_DEC_ERR_Q0_0_INTRO_175_err_intro_q0_0_175(o_LDPC_DEC_ERR_Q0_0_INTRO_175_err_intro_q0_0_175),
.o_LDPC_DEC_ERR_Q0_0_INTRO_176_err_intro_q0_0_176(o_LDPC_DEC_ERR_Q0_0_INTRO_176_err_intro_q0_0_176),
.o_LDPC_DEC_ERR_Q0_0_INTRO_177_err_intro_q0_0_177(o_LDPC_DEC_ERR_Q0_0_INTRO_177_err_intro_q0_0_177),
.o_LDPC_DEC_ERR_Q0_0_INTRO_178_err_intro_q0_0_178(o_LDPC_DEC_ERR_Q0_0_INTRO_178_err_intro_q0_0_178),
.o_LDPC_DEC_ERR_Q0_0_INTRO_179_err_intro_q0_0_179(o_LDPC_DEC_ERR_Q0_0_INTRO_179_err_intro_q0_0_179),
.o_LDPC_DEC_ERR_Q0_0_INTRO_180_err_intro_q0_0_180(o_LDPC_DEC_ERR_Q0_0_INTRO_180_err_intro_q0_0_180),
.o_LDPC_DEC_ERR_Q0_0_INTRO_181_err_intro_q0_0_181(o_LDPC_DEC_ERR_Q0_0_INTRO_181_err_intro_q0_0_181),
.o_LDPC_DEC_ERR_Q0_0_INTRO_182_err_intro_q0_0_182(o_LDPC_DEC_ERR_Q0_0_INTRO_182_err_intro_q0_0_182),
.o_LDPC_DEC_ERR_Q0_0_INTRO_183_err_intro_q0_0_183(o_LDPC_DEC_ERR_Q0_0_INTRO_183_err_intro_q0_0_183),
.o_LDPC_DEC_ERR_Q0_0_INTRO_184_err_intro_q0_0_184(o_LDPC_DEC_ERR_Q0_0_INTRO_184_err_intro_q0_0_184),
.o_LDPC_DEC_ERR_Q0_0_INTRO_185_err_intro_q0_0_185(o_LDPC_DEC_ERR_Q0_0_INTRO_185_err_intro_q0_0_185),
.o_LDPC_DEC_ERR_Q0_0_INTRO_186_err_intro_q0_0_186(o_LDPC_DEC_ERR_Q0_0_INTRO_186_err_intro_q0_0_186),
.o_LDPC_DEC_ERR_Q0_0_INTRO_187_err_intro_q0_0_187(o_LDPC_DEC_ERR_Q0_0_INTRO_187_err_intro_q0_0_187),
.o_LDPC_DEC_ERR_Q0_0_INTRO_188_err_intro_q0_0_188(o_LDPC_DEC_ERR_Q0_0_INTRO_188_err_intro_q0_0_188),
.o_LDPC_DEC_ERR_Q0_0_INTRO_189_err_intro_q0_0_189(o_LDPC_DEC_ERR_Q0_0_INTRO_189_err_intro_q0_0_189),
.o_LDPC_DEC_ERR_Q0_0_INTRO_190_err_intro_q0_0_190(o_LDPC_DEC_ERR_Q0_0_INTRO_190_err_intro_q0_0_190),
.o_LDPC_DEC_ERR_Q0_0_INTRO_191_err_intro_q0_0_191(o_LDPC_DEC_ERR_Q0_0_INTRO_191_err_intro_q0_0_191),
.o_LDPC_DEC_ERR_Q0_0_INTRO_192_err_intro_q0_0_192(o_LDPC_DEC_ERR_Q0_0_INTRO_192_err_intro_q0_0_192),
.o_LDPC_DEC_ERR_Q0_0_INTRO_193_err_intro_q0_0_193(o_LDPC_DEC_ERR_Q0_0_INTRO_193_err_intro_q0_0_193),
.o_LDPC_DEC_ERR_Q0_0_INTRO_194_err_intro_q0_0_194(o_LDPC_DEC_ERR_Q0_0_INTRO_194_err_intro_q0_0_194),
.o_LDPC_DEC_ERR_Q0_0_INTRO_195_err_intro_q0_0_195(o_LDPC_DEC_ERR_Q0_0_INTRO_195_err_intro_q0_0_195),
.o_LDPC_DEC_ERR_Q0_0_INTRO_196_err_intro_q0_0_196(o_LDPC_DEC_ERR_Q0_0_INTRO_196_err_intro_q0_0_196),
.o_LDPC_DEC_ERR_Q0_0_INTRO_197_err_intro_q0_0_197(o_LDPC_DEC_ERR_Q0_0_INTRO_197_err_intro_q0_0_197),
.o_LDPC_DEC_ERR_Q0_0_INTRO_198_err_intro_q0_0_198(o_LDPC_DEC_ERR_Q0_0_INTRO_198_err_intro_q0_0_198),
.o_LDPC_DEC_ERR_Q0_0_INTRO_199_err_intro_q0_0_199(o_LDPC_DEC_ERR_Q0_0_INTRO_199_err_intro_q0_0_199),
.o_LDPC_DEC_ERR_Q0_0_INTRO_200_err_intro_q0_0_200(o_LDPC_DEC_ERR_Q0_0_INTRO_200_err_intro_q0_0_200),
.o_LDPC_DEC_ERR_Q0_0_INTRO_201_err_intro_q0_0_201(o_LDPC_DEC_ERR_Q0_0_INTRO_201_err_intro_q0_0_201),
.o_LDPC_DEC_ERR_Q0_0_INTRO_202_err_intro_q0_0_202(o_LDPC_DEC_ERR_Q0_0_INTRO_202_err_intro_q0_0_202),
.o_LDPC_DEC_ERR_Q0_0_INTRO_203_err_intro_q0_0_203(o_LDPC_DEC_ERR_Q0_0_INTRO_203_err_intro_q0_0_203),
.o_LDPC_DEC_ERR_Q0_0_INTRO_204_err_intro_q0_0_204(o_LDPC_DEC_ERR_Q0_0_INTRO_204_err_intro_q0_0_204),
.o_LDPC_DEC_ERR_Q0_0_INTRO_205_err_intro_q0_0_205(o_LDPC_DEC_ERR_Q0_0_INTRO_205_err_intro_q0_0_205),
.o_LDPC_DEC_ERR_Q0_0_INTRO_206_err_intro_q0_0_206(o_LDPC_DEC_ERR_Q0_0_INTRO_206_err_intro_q0_0_206),
.o_LDPC_DEC_ERR_Q0_0_INTRO_207_err_intro_q0_0_207(o_LDPC_DEC_ERR_Q0_0_INTRO_207_err_intro_q0_0_207),
.o_LDPC_DEC_ERR_Q0_1_INTRO_0_err_intro_q0_1_0(o_LDPC_DEC_ERR_Q0_1_INTRO_0_err_intro_q0_1_0),
.o_LDPC_DEC_ERR_Q0_1_INTRO_1_err_intro_q0_1_1(o_LDPC_DEC_ERR_Q0_1_INTRO_1_err_intro_q0_1_1),
.o_LDPC_DEC_ERR_Q0_1_INTRO_2_err_intro_q0_1_2(o_LDPC_DEC_ERR_Q0_1_INTRO_2_err_intro_q0_1_2),
.o_LDPC_DEC_ERR_Q0_1_INTRO_3_err_intro_q0_1_3(o_LDPC_DEC_ERR_Q0_1_INTRO_3_err_intro_q0_1_3),
.o_LDPC_DEC_ERR_Q0_1_INTRO_4_err_intro_q0_1_4(o_LDPC_DEC_ERR_Q0_1_INTRO_4_err_intro_q0_1_4),
.o_LDPC_DEC_ERR_Q0_1_INTRO_5_err_intro_q0_1_5(o_LDPC_DEC_ERR_Q0_1_INTRO_5_err_intro_q0_1_5),
.o_LDPC_DEC_ERR_Q0_1_INTRO_6_err_intro_q0_1_6(o_LDPC_DEC_ERR_Q0_1_INTRO_6_err_intro_q0_1_6),
.o_LDPC_DEC_ERR_Q0_1_INTRO_7_err_intro_q0_1_7(o_LDPC_DEC_ERR_Q0_1_INTRO_7_err_intro_q0_1_7),
.o_LDPC_DEC_ERR_Q0_1_INTRO_8_err_intro_q0_1_8(o_LDPC_DEC_ERR_Q0_1_INTRO_8_err_intro_q0_1_8),
.o_LDPC_DEC_ERR_Q0_1_INTRO_9_err_intro_q0_1_9(o_LDPC_DEC_ERR_Q0_1_INTRO_9_err_intro_q0_1_9),
.o_LDPC_DEC_ERR_Q0_1_INTRO_10_err_intro_q0_1_10(o_LDPC_DEC_ERR_Q0_1_INTRO_10_err_intro_q0_1_10),
.o_LDPC_DEC_ERR_Q0_1_INTRO_11_err_intro_q0_1_11(o_LDPC_DEC_ERR_Q0_1_INTRO_11_err_intro_q0_1_11),
.o_LDPC_DEC_ERR_Q0_1_INTRO_12_err_intro_q0_1_12(o_LDPC_DEC_ERR_Q0_1_INTRO_12_err_intro_q0_1_12),
.o_LDPC_DEC_ERR_Q0_1_INTRO_13_err_intro_q0_1_13(o_LDPC_DEC_ERR_Q0_1_INTRO_13_err_intro_q0_1_13),
.o_LDPC_DEC_ERR_Q0_1_INTRO_14_err_intro_q0_1_14(o_LDPC_DEC_ERR_Q0_1_INTRO_14_err_intro_q0_1_14),
.o_LDPC_DEC_ERR_Q0_1_INTRO_15_err_intro_q0_1_15(o_LDPC_DEC_ERR_Q0_1_INTRO_15_err_intro_q0_1_15),
.o_LDPC_DEC_ERR_Q0_1_INTRO_16_err_intro_q0_1_16(o_LDPC_DEC_ERR_Q0_1_INTRO_16_err_intro_q0_1_16),
.o_LDPC_DEC_ERR_Q0_1_INTRO_17_err_intro_q0_1_17(o_LDPC_DEC_ERR_Q0_1_INTRO_17_err_intro_q0_1_17),
.o_LDPC_DEC_ERR_Q0_1_INTRO_18_err_intro_q0_1_18(o_LDPC_DEC_ERR_Q0_1_INTRO_18_err_intro_q0_1_18),
.o_LDPC_DEC_ERR_Q0_1_INTRO_19_err_intro_q0_1_19(o_LDPC_DEC_ERR_Q0_1_INTRO_19_err_intro_q0_1_19),
.o_LDPC_DEC_ERR_Q0_1_INTRO_20_err_intro_q0_1_20(o_LDPC_DEC_ERR_Q0_1_INTRO_20_err_intro_q0_1_20),
.o_LDPC_DEC_ERR_Q0_1_INTRO_21_err_intro_q0_1_21(o_LDPC_DEC_ERR_Q0_1_INTRO_21_err_intro_q0_1_21),
.o_LDPC_DEC_ERR_Q0_1_INTRO_22_err_intro_q0_1_22(o_LDPC_DEC_ERR_Q0_1_INTRO_22_err_intro_q0_1_22),
.o_LDPC_DEC_ERR_Q0_1_INTRO_23_err_intro_q0_1_23(o_LDPC_DEC_ERR_Q0_1_INTRO_23_err_intro_q0_1_23),
.o_LDPC_DEC_ERR_Q0_1_INTRO_24_err_intro_q0_1_24(o_LDPC_DEC_ERR_Q0_1_INTRO_24_err_intro_q0_1_24),
.o_LDPC_DEC_ERR_Q0_1_INTRO_25_err_intro_q0_1_25(o_LDPC_DEC_ERR_Q0_1_INTRO_25_err_intro_q0_1_25),
.o_LDPC_DEC_ERR_Q0_1_INTRO_26_err_intro_q0_1_26(o_LDPC_DEC_ERR_Q0_1_INTRO_26_err_intro_q0_1_26),
.o_LDPC_DEC_ERR_Q0_1_INTRO_27_err_intro_q0_1_27(o_LDPC_DEC_ERR_Q0_1_INTRO_27_err_intro_q0_1_27),
.o_LDPC_DEC_ERR_Q0_1_INTRO_28_err_intro_q0_1_28(o_LDPC_DEC_ERR_Q0_1_INTRO_28_err_intro_q0_1_28),
.o_LDPC_DEC_ERR_Q0_1_INTRO_29_err_intro_q0_1_29(o_LDPC_DEC_ERR_Q0_1_INTRO_29_err_intro_q0_1_29),
.o_LDPC_DEC_ERR_Q0_1_INTRO_30_err_intro_q0_1_30(o_LDPC_DEC_ERR_Q0_1_INTRO_30_err_intro_q0_1_30),
.o_LDPC_DEC_ERR_Q0_1_INTRO_31_err_intro_q0_1_31(o_LDPC_DEC_ERR_Q0_1_INTRO_31_err_intro_q0_1_31),
.o_LDPC_DEC_ERR_Q0_1_INTRO_32_err_intro_q0_1_32(o_LDPC_DEC_ERR_Q0_1_INTRO_32_err_intro_q0_1_32),
.o_LDPC_DEC_ERR_Q0_1_INTRO_33_err_intro_q0_1_33(o_LDPC_DEC_ERR_Q0_1_INTRO_33_err_intro_q0_1_33),
.o_LDPC_DEC_ERR_Q0_1_INTRO_34_err_intro_q0_1_34(o_LDPC_DEC_ERR_Q0_1_INTRO_34_err_intro_q0_1_34),
.o_LDPC_DEC_ERR_Q0_1_INTRO_35_err_intro_q0_1_35(o_LDPC_DEC_ERR_Q0_1_INTRO_35_err_intro_q0_1_35),
.o_LDPC_DEC_ERR_Q0_1_INTRO_36_err_intro_q0_1_36(o_LDPC_DEC_ERR_Q0_1_INTRO_36_err_intro_q0_1_36),
.o_LDPC_DEC_ERR_Q0_1_INTRO_37_err_intro_q0_1_37(o_LDPC_DEC_ERR_Q0_1_INTRO_37_err_intro_q0_1_37),
.o_LDPC_DEC_ERR_Q0_1_INTRO_38_err_intro_q0_1_38(o_LDPC_DEC_ERR_Q0_1_INTRO_38_err_intro_q0_1_38),
.o_LDPC_DEC_ERR_Q0_1_INTRO_39_err_intro_q0_1_39(o_LDPC_DEC_ERR_Q0_1_INTRO_39_err_intro_q0_1_39),
.o_LDPC_DEC_ERR_Q0_1_INTRO_40_err_intro_q0_1_40(o_LDPC_DEC_ERR_Q0_1_INTRO_40_err_intro_q0_1_40),
.o_LDPC_DEC_ERR_Q0_1_INTRO_41_err_intro_q0_1_41(o_LDPC_DEC_ERR_Q0_1_INTRO_41_err_intro_q0_1_41),
.o_LDPC_DEC_ERR_Q0_1_INTRO_42_err_intro_q0_1_42(o_LDPC_DEC_ERR_Q0_1_INTRO_42_err_intro_q0_1_42),
.o_LDPC_DEC_ERR_Q0_1_INTRO_43_err_intro_q0_1_43(o_LDPC_DEC_ERR_Q0_1_INTRO_43_err_intro_q0_1_43),
.o_LDPC_DEC_ERR_Q0_1_INTRO_44_err_intro_q0_1_44(o_LDPC_DEC_ERR_Q0_1_INTRO_44_err_intro_q0_1_44),
.o_LDPC_DEC_ERR_Q0_1_INTRO_45_err_intro_q0_1_45(o_LDPC_DEC_ERR_Q0_1_INTRO_45_err_intro_q0_1_45),
.o_LDPC_DEC_ERR_Q0_1_INTRO_46_err_intro_q0_1_46(o_LDPC_DEC_ERR_Q0_1_INTRO_46_err_intro_q0_1_46),
.o_LDPC_DEC_ERR_Q0_1_INTRO_47_err_intro_q0_1_47(o_LDPC_DEC_ERR_Q0_1_INTRO_47_err_intro_q0_1_47),
.o_LDPC_DEC_ERR_Q0_1_INTRO_48_err_intro_q0_1_48(o_LDPC_DEC_ERR_Q0_1_INTRO_48_err_intro_q0_1_48),
.o_LDPC_DEC_ERR_Q0_1_INTRO_49_err_intro_q0_1_49(o_LDPC_DEC_ERR_Q0_1_INTRO_49_err_intro_q0_1_49),
.o_LDPC_DEC_ERR_Q0_1_INTRO_50_err_intro_q0_1_50(o_LDPC_DEC_ERR_Q0_1_INTRO_50_err_intro_q0_1_50),
.o_LDPC_DEC_ERR_Q0_1_INTRO_51_err_intro_q0_1_51(o_LDPC_DEC_ERR_Q0_1_INTRO_51_err_intro_q0_1_51),
.o_LDPC_DEC_ERR_Q0_1_INTRO_52_err_intro_q0_1_52(o_LDPC_DEC_ERR_Q0_1_INTRO_52_err_intro_q0_1_52),
.o_LDPC_DEC_ERR_Q0_1_INTRO_53_err_intro_q0_1_53(o_LDPC_DEC_ERR_Q0_1_INTRO_53_err_intro_q0_1_53),
.o_LDPC_DEC_ERR_Q0_1_INTRO_54_err_intro_q0_1_54(o_LDPC_DEC_ERR_Q0_1_INTRO_54_err_intro_q0_1_54),
.o_LDPC_DEC_ERR_Q0_1_INTRO_55_err_intro_q0_1_55(o_LDPC_DEC_ERR_Q0_1_INTRO_55_err_intro_q0_1_55),
.o_LDPC_DEC_ERR_Q0_1_INTRO_56_err_intro_q0_1_56(o_LDPC_DEC_ERR_Q0_1_INTRO_56_err_intro_q0_1_56),
.o_LDPC_DEC_ERR_Q0_1_INTRO_57_err_intro_q0_1_57(o_LDPC_DEC_ERR_Q0_1_INTRO_57_err_intro_q0_1_57),
.o_LDPC_DEC_ERR_Q0_1_INTRO_58_err_intro_q0_1_58(o_LDPC_DEC_ERR_Q0_1_INTRO_58_err_intro_q0_1_58),
.o_LDPC_DEC_ERR_Q0_1_INTRO_59_err_intro_q0_1_59(o_LDPC_DEC_ERR_Q0_1_INTRO_59_err_intro_q0_1_59),
.o_LDPC_DEC_ERR_Q0_1_INTRO_60_err_intro_q0_1_60(o_LDPC_DEC_ERR_Q0_1_INTRO_60_err_intro_q0_1_60),
.o_LDPC_DEC_ERR_Q0_1_INTRO_61_err_intro_q0_1_61(o_LDPC_DEC_ERR_Q0_1_INTRO_61_err_intro_q0_1_61),
.o_LDPC_DEC_ERR_Q0_1_INTRO_62_err_intro_q0_1_62(o_LDPC_DEC_ERR_Q0_1_INTRO_62_err_intro_q0_1_62),
.o_LDPC_DEC_ERR_Q0_1_INTRO_63_err_intro_q0_1_63(o_LDPC_DEC_ERR_Q0_1_INTRO_63_err_intro_q0_1_63),
.o_LDPC_DEC_ERR_Q0_1_INTRO_64_err_intro_q0_1_64(o_LDPC_DEC_ERR_Q0_1_INTRO_64_err_intro_q0_1_64),
.o_LDPC_DEC_ERR_Q0_1_INTRO_65_err_intro_q0_1_65(o_LDPC_DEC_ERR_Q0_1_INTRO_65_err_intro_q0_1_65),
.o_LDPC_DEC_ERR_Q0_1_INTRO_66_err_intro_q0_1_66(o_LDPC_DEC_ERR_Q0_1_INTRO_66_err_intro_q0_1_66),
.o_LDPC_DEC_ERR_Q0_1_INTRO_67_err_intro_q0_1_67(o_LDPC_DEC_ERR_Q0_1_INTRO_67_err_intro_q0_1_67),
.o_LDPC_DEC_ERR_Q0_1_INTRO_68_err_intro_q0_1_68(o_LDPC_DEC_ERR_Q0_1_INTRO_68_err_intro_q0_1_68),
.o_LDPC_DEC_ERR_Q0_1_INTRO_69_err_intro_q0_1_69(o_LDPC_DEC_ERR_Q0_1_INTRO_69_err_intro_q0_1_69),
.o_LDPC_DEC_ERR_Q0_1_INTRO_70_err_intro_q0_1_70(o_LDPC_DEC_ERR_Q0_1_INTRO_70_err_intro_q0_1_70),
.o_LDPC_DEC_ERR_Q0_1_INTRO_71_err_intro_q0_1_71(o_LDPC_DEC_ERR_Q0_1_INTRO_71_err_intro_q0_1_71),
.o_LDPC_DEC_ERR_Q0_1_INTRO_72_err_intro_q0_1_72(o_LDPC_DEC_ERR_Q0_1_INTRO_72_err_intro_q0_1_72),
.o_LDPC_DEC_ERR_Q0_1_INTRO_73_err_intro_q0_1_73(o_LDPC_DEC_ERR_Q0_1_INTRO_73_err_intro_q0_1_73),
.o_LDPC_DEC_ERR_Q0_1_INTRO_74_err_intro_q0_1_74(o_LDPC_DEC_ERR_Q0_1_INTRO_74_err_intro_q0_1_74),
.o_LDPC_DEC_ERR_Q0_1_INTRO_75_err_intro_q0_1_75(o_LDPC_DEC_ERR_Q0_1_INTRO_75_err_intro_q0_1_75),
.o_LDPC_DEC_ERR_Q0_1_INTRO_76_err_intro_q0_1_76(o_LDPC_DEC_ERR_Q0_1_INTRO_76_err_intro_q0_1_76),
.o_LDPC_DEC_ERR_Q0_1_INTRO_77_err_intro_q0_1_77(o_LDPC_DEC_ERR_Q0_1_INTRO_77_err_intro_q0_1_77),
.o_LDPC_DEC_ERR_Q0_1_INTRO_78_err_intro_q0_1_78(o_LDPC_DEC_ERR_Q0_1_INTRO_78_err_intro_q0_1_78),
.o_LDPC_DEC_ERR_Q0_1_INTRO_79_err_intro_q0_1_79(o_LDPC_DEC_ERR_Q0_1_INTRO_79_err_intro_q0_1_79),
.o_LDPC_DEC_ERR_Q0_1_INTRO_80_err_intro_q0_1_80(o_LDPC_DEC_ERR_Q0_1_INTRO_80_err_intro_q0_1_80),
.o_LDPC_DEC_ERR_Q0_1_INTRO_81_err_intro_q0_1_81(o_LDPC_DEC_ERR_Q0_1_INTRO_81_err_intro_q0_1_81),
.o_LDPC_DEC_ERR_Q0_1_INTRO_82_err_intro_q0_1_82(o_LDPC_DEC_ERR_Q0_1_INTRO_82_err_intro_q0_1_82),
.o_LDPC_DEC_ERR_Q0_1_INTRO_83_err_intro_q0_1_83(o_LDPC_DEC_ERR_Q0_1_INTRO_83_err_intro_q0_1_83),
.o_LDPC_DEC_ERR_Q0_1_INTRO_84_err_intro_q0_1_84(o_LDPC_DEC_ERR_Q0_1_INTRO_84_err_intro_q0_1_84),
.o_LDPC_DEC_ERR_Q0_1_INTRO_85_err_intro_q0_1_85(o_LDPC_DEC_ERR_Q0_1_INTRO_85_err_intro_q0_1_85),
.o_LDPC_DEC_ERR_Q0_1_INTRO_86_err_intro_q0_1_86(o_LDPC_DEC_ERR_Q0_1_INTRO_86_err_intro_q0_1_86),
.o_LDPC_DEC_ERR_Q0_1_INTRO_87_err_intro_q0_1_87(o_LDPC_DEC_ERR_Q0_1_INTRO_87_err_intro_q0_1_87),
.o_LDPC_DEC_ERR_Q0_1_INTRO_88_err_intro_q0_1_88(o_LDPC_DEC_ERR_Q0_1_INTRO_88_err_intro_q0_1_88),
.o_LDPC_DEC_ERR_Q0_1_INTRO_89_err_intro_q0_1_89(o_LDPC_DEC_ERR_Q0_1_INTRO_89_err_intro_q0_1_89),
.o_LDPC_DEC_ERR_Q0_1_INTRO_90_err_intro_q0_1_90(o_LDPC_DEC_ERR_Q0_1_INTRO_90_err_intro_q0_1_90),
.o_LDPC_DEC_ERR_Q0_1_INTRO_91_err_intro_q0_1_91(o_LDPC_DEC_ERR_Q0_1_INTRO_91_err_intro_q0_1_91),
.o_LDPC_DEC_ERR_Q0_1_INTRO_92_err_intro_q0_1_92(o_LDPC_DEC_ERR_Q0_1_INTRO_92_err_intro_q0_1_92),
.o_LDPC_DEC_ERR_Q0_1_INTRO_93_err_intro_q0_1_93(o_LDPC_DEC_ERR_Q0_1_INTRO_93_err_intro_q0_1_93),
.o_LDPC_DEC_ERR_Q0_1_INTRO_94_err_intro_q0_1_94(o_LDPC_DEC_ERR_Q0_1_INTRO_94_err_intro_q0_1_94),
.o_LDPC_DEC_ERR_Q0_1_INTRO_95_err_intro_q0_1_95(o_LDPC_DEC_ERR_Q0_1_INTRO_95_err_intro_q0_1_95),
.o_LDPC_DEC_ERR_Q0_1_INTRO_96_err_intro_q0_1_96(o_LDPC_DEC_ERR_Q0_1_INTRO_96_err_intro_q0_1_96),
.o_LDPC_DEC_ERR_Q0_1_INTRO_97_err_intro_q0_1_97(o_LDPC_DEC_ERR_Q0_1_INTRO_97_err_intro_q0_1_97),
.o_LDPC_DEC_ERR_Q0_1_INTRO_98_err_intro_q0_1_98(o_LDPC_DEC_ERR_Q0_1_INTRO_98_err_intro_q0_1_98),
.o_LDPC_DEC_ERR_Q0_1_INTRO_99_err_intro_q0_1_99(o_LDPC_DEC_ERR_Q0_1_INTRO_99_err_intro_q0_1_99),
.o_LDPC_DEC_ERR_Q0_1_INTRO_100_err_intro_q0_1_100(o_LDPC_DEC_ERR_Q0_1_INTRO_100_err_intro_q0_1_100),
.o_LDPC_DEC_ERR_Q0_1_INTRO_101_err_intro_q0_1_101(o_LDPC_DEC_ERR_Q0_1_INTRO_101_err_intro_q0_1_101),
.o_LDPC_DEC_ERR_Q0_1_INTRO_102_err_intro_q0_1_102(o_LDPC_DEC_ERR_Q0_1_INTRO_102_err_intro_q0_1_102),
.o_LDPC_DEC_ERR_Q0_1_INTRO_103_err_intro_q0_1_103(o_LDPC_DEC_ERR_Q0_1_INTRO_103_err_intro_q0_1_103),
.o_LDPC_DEC_ERR_Q0_1_INTRO_104_err_intro_q0_1_104(o_LDPC_DEC_ERR_Q0_1_INTRO_104_err_intro_q0_1_104),
.o_LDPC_DEC_ERR_Q0_1_INTRO_105_err_intro_q0_1_105(o_LDPC_DEC_ERR_Q0_1_INTRO_105_err_intro_q0_1_105),
.o_LDPC_DEC_ERR_Q0_1_INTRO_106_err_intro_q0_1_106(o_LDPC_DEC_ERR_Q0_1_INTRO_106_err_intro_q0_1_106),
.o_LDPC_DEC_ERR_Q0_1_INTRO_107_err_intro_q0_1_107(o_LDPC_DEC_ERR_Q0_1_INTRO_107_err_intro_q0_1_107),
.o_LDPC_DEC_ERR_Q0_1_INTRO_108_err_intro_q0_1_108(o_LDPC_DEC_ERR_Q0_1_INTRO_108_err_intro_q0_1_108),
.o_LDPC_DEC_ERR_Q0_1_INTRO_109_err_intro_q0_1_109(o_LDPC_DEC_ERR_Q0_1_INTRO_109_err_intro_q0_1_109),
.o_LDPC_DEC_ERR_Q0_1_INTRO_110_err_intro_q0_1_110(o_LDPC_DEC_ERR_Q0_1_INTRO_110_err_intro_q0_1_110),
.o_LDPC_DEC_ERR_Q0_1_INTRO_111_err_intro_q0_1_111(o_LDPC_DEC_ERR_Q0_1_INTRO_111_err_intro_q0_1_111),
.o_LDPC_DEC_ERR_Q0_1_INTRO_112_err_intro_q0_1_112(o_LDPC_DEC_ERR_Q0_1_INTRO_112_err_intro_q0_1_112),
.o_LDPC_DEC_ERR_Q0_1_INTRO_113_err_intro_q0_1_113(o_LDPC_DEC_ERR_Q0_1_INTRO_113_err_intro_q0_1_113),
.o_LDPC_DEC_ERR_Q0_1_INTRO_114_err_intro_q0_1_114(o_LDPC_DEC_ERR_Q0_1_INTRO_114_err_intro_q0_1_114),
.o_LDPC_DEC_ERR_Q0_1_INTRO_115_err_intro_q0_1_115(o_LDPC_DEC_ERR_Q0_1_INTRO_115_err_intro_q0_1_115),
.o_LDPC_DEC_ERR_Q0_1_INTRO_116_err_intro_q0_1_116(o_LDPC_DEC_ERR_Q0_1_INTRO_116_err_intro_q0_1_116),
.o_LDPC_DEC_ERR_Q0_1_INTRO_117_err_intro_q0_1_117(o_LDPC_DEC_ERR_Q0_1_INTRO_117_err_intro_q0_1_117),
.o_LDPC_DEC_ERR_Q0_1_INTRO_118_err_intro_q0_1_118(o_LDPC_DEC_ERR_Q0_1_INTRO_118_err_intro_q0_1_118),
.o_LDPC_DEC_ERR_Q0_1_INTRO_119_err_intro_q0_1_119(o_LDPC_DEC_ERR_Q0_1_INTRO_119_err_intro_q0_1_119),
.o_LDPC_DEC_ERR_Q0_1_INTRO_120_err_intro_q0_1_120(o_LDPC_DEC_ERR_Q0_1_INTRO_120_err_intro_q0_1_120),
.o_LDPC_DEC_ERR_Q0_1_INTRO_121_err_intro_q0_1_121(o_LDPC_DEC_ERR_Q0_1_INTRO_121_err_intro_q0_1_121),
.o_LDPC_DEC_ERR_Q0_1_INTRO_122_err_intro_q0_1_122(o_LDPC_DEC_ERR_Q0_1_INTRO_122_err_intro_q0_1_122),
.o_LDPC_DEC_ERR_Q0_1_INTRO_123_err_intro_q0_1_123(o_LDPC_DEC_ERR_Q0_1_INTRO_123_err_intro_q0_1_123),
.o_LDPC_DEC_ERR_Q0_1_INTRO_124_err_intro_q0_1_124(o_LDPC_DEC_ERR_Q0_1_INTRO_124_err_intro_q0_1_124),
.o_LDPC_DEC_ERR_Q0_1_INTRO_125_err_intro_q0_1_125(o_LDPC_DEC_ERR_Q0_1_INTRO_125_err_intro_q0_1_125),
.o_LDPC_DEC_ERR_Q0_1_INTRO_126_err_intro_q0_1_126(o_LDPC_DEC_ERR_Q0_1_INTRO_126_err_intro_q0_1_126),
.o_LDPC_DEC_ERR_Q0_1_INTRO_127_err_intro_q0_1_127(o_LDPC_DEC_ERR_Q0_1_INTRO_127_err_intro_q0_1_127),
.o_LDPC_DEC_ERR_Q0_1_INTRO_128_err_intro_q0_1_128(o_LDPC_DEC_ERR_Q0_1_INTRO_128_err_intro_q0_1_128),
.o_LDPC_DEC_ERR_Q0_1_INTRO_129_err_intro_q0_1_129(o_LDPC_DEC_ERR_Q0_1_INTRO_129_err_intro_q0_1_129),
.o_LDPC_DEC_ERR_Q0_1_INTRO_130_err_intro_q0_1_130(o_LDPC_DEC_ERR_Q0_1_INTRO_130_err_intro_q0_1_130),
.o_LDPC_DEC_ERR_Q0_1_INTRO_131_err_intro_q0_1_131(o_LDPC_DEC_ERR_Q0_1_INTRO_131_err_intro_q0_1_131),
.o_LDPC_DEC_ERR_Q0_1_INTRO_132_err_intro_q0_1_132(o_LDPC_DEC_ERR_Q0_1_INTRO_132_err_intro_q0_1_132),
.o_LDPC_DEC_ERR_Q0_1_INTRO_133_err_intro_q0_1_133(o_LDPC_DEC_ERR_Q0_1_INTRO_133_err_intro_q0_1_133),
.o_LDPC_DEC_ERR_Q0_1_INTRO_134_err_intro_q0_1_134(o_LDPC_DEC_ERR_Q0_1_INTRO_134_err_intro_q0_1_134),
.o_LDPC_DEC_ERR_Q0_1_INTRO_135_err_intro_q0_1_135(o_LDPC_DEC_ERR_Q0_1_INTRO_135_err_intro_q0_1_135),
.o_LDPC_DEC_ERR_Q0_1_INTRO_136_err_intro_q0_1_136(o_LDPC_DEC_ERR_Q0_1_INTRO_136_err_intro_q0_1_136),
.o_LDPC_DEC_ERR_Q0_1_INTRO_137_err_intro_q0_1_137(o_LDPC_DEC_ERR_Q0_1_INTRO_137_err_intro_q0_1_137),
.o_LDPC_DEC_ERR_Q0_1_INTRO_138_err_intro_q0_1_138(o_LDPC_DEC_ERR_Q0_1_INTRO_138_err_intro_q0_1_138),
.o_LDPC_DEC_ERR_Q0_1_INTRO_139_err_intro_q0_1_139(o_LDPC_DEC_ERR_Q0_1_INTRO_139_err_intro_q0_1_139),
.o_LDPC_DEC_ERR_Q0_1_INTRO_140_err_intro_q0_1_140(o_LDPC_DEC_ERR_Q0_1_INTRO_140_err_intro_q0_1_140),
.o_LDPC_DEC_ERR_Q0_1_INTRO_141_err_intro_q0_1_141(o_LDPC_DEC_ERR_Q0_1_INTRO_141_err_intro_q0_1_141),
.o_LDPC_DEC_ERR_Q0_1_INTRO_142_err_intro_q0_1_142(o_LDPC_DEC_ERR_Q0_1_INTRO_142_err_intro_q0_1_142),
.o_LDPC_DEC_ERR_Q0_1_INTRO_143_err_intro_q0_1_143(o_LDPC_DEC_ERR_Q0_1_INTRO_143_err_intro_q0_1_143),
.o_LDPC_DEC_ERR_Q0_1_INTRO_144_err_intro_q0_1_144(o_LDPC_DEC_ERR_Q0_1_INTRO_144_err_intro_q0_1_144),
.o_LDPC_DEC_ERR_Q0_1_INTRO_145_err_intro_q0_1_145(o_LDPC_DEC_ERR_Q0_1_INTRO_145_err_intro_q0_1_145),
.o_LDPC_DEC_ERR_Q0_1_INTRO_146_err_intro_q0_1_146(o_LDPC_DEC_ERR_Q0_1_INTRO_146_err_intro_q0_1_146),
.o_LDPC_DEC_ERR_Q0_1_INTRO_147_err_intro_q0_1_147(o_LDPC_DEC_ERR_Q0_1_INTRO_147_err_intro_q0_1_147),
.o_LDPC_DEC_ERR_Q0_1_INTRO_148_err_intro_q0_1_148(o_LDPC_DEC_ERR_Q0_1_INTRO_148_err_intro_q0_1_148),
.o_LDPC_DEC_ERR_Q0_1_INTRO_149_err_intro_q0_1_149(o_LDPC_DEC_ERR_Q0_1_INTRO_149_err_intro_q0_1_149),
.o_LDPC_DEC_ERR_Q0_1_INTRO_150_err_intro_q0_1_150(o_LDPC_DEC_ERR_Q0_1_INTRO_150_err_intro_q0_1_150),
.o_LDPC_DEC_ERR_Q0_1_INTRO_151_err_intro_q0_1_151(o_LDPC_DEC_ERR_Q0_1_INTRO_151_err_intro_q0_1_151),
.o_LDPC_DEC_ERR_Q0_1_INTRO_152_err_intro_q0_1_152(o_LDPC_DEC_ERR_Q0_1_INTRO_152_err_intro_q0_1_152),
.o_LDPC_DEC_ERR_Q0_1_INTRO_153_err_intro_q0_1_153(o_LDPC_DEC_ERR_Q0_1_INTRO_153_err_intro_q0_1_153),
.o_LDPC_DEC_ERR_Q0_1_INTRO_154_err_intro_q0_1_154(o_LDPC_DEC_ERR_Q0_1_INTRO_154_err_intro_q0_1_154),
.o_LDPC_DEC_ERR_Q0_1_INTRO_155_err_intro_q0_1_155(o_LDPC_DEC_ERR_Q0_1_INTRO_155_err_intro_q0_1_155),
.o_LDPC_DEC_ERR_Q0_1_INTRO_156_err_intro_q0_1_156(o_LDPC_DEC_ERR_Q0_1_INTRO_156_err_intro_q0_1_156),
.o_LDPC_DEC_ERR_Q0_1_INTRO_157_err_intro_q0_1_157(o_LDPC_DEC_ERR_Q0_1_INTRO_157_err_intro_q0_1_157),
.o_LDPC_DEC_ERR_Q0_1_INTRO_158_err_intro_q0_1_158(o_LDPC_DEC_ERR_Q0_1_INTRO_158_err_intro_q0_1_158),
.o_LDPC_DEC_ERR_Q0_1_INTRO_159_err_intro_q0_1_159(o_LDPC_DEC_ERR_Q0_1_INTRO_159_err_intro_q0_1_159),
.o_LDPC_DEC_ERR_Q0_1_INTRO_160_err_intro_q0_1_160(o_LDPC_DEC_ERR_Q0_1_INTRO_160_err_intro_q0_1_160),
.o_LDPC_DEC_ERR_Q0_1_INTRO_161_err_intro_q0_1_161(o_LDPC_DEC_ERR_Q0_1_INTRO_161_err_intro_q0_1_161),
.o_LDPC_DEC_ERR_Q0_1_INTRO_162_err_intro_q0_1_162(o_LDPC_DEC_ERR_Q0_1_INTRO_162_err_intro_q0_1_162),
.o_LDPC_DEC_ERR_Q0_1_INTRO_163_err_intro_q0_1_163(o_LDPC_DEC_ERR_Q0_1_INTRO_163_err_intro_q0_1_163),
.o_LDPC_DEC_ERR_Q0_1_INTRO_164_err_intro_q0_1_164(o_LDPC_DEC_ERR_Q0_1_INTRO_164_err_intro_q0_1_164),
.o_LDPC_DEC_ERR_Q0_1_INTRO_165_err_intro_q0_1_165(o_LDPC_DEC_ERR_Q0_1_INTRO_165_err_intro_q0_1_165),
.o_LDPC_DEC_ERR_Q0_1_INTRO_166_err_intro_q0_1_166(o_LDPC_DEC_ERR_Q0_1_INTRO_166_err_intro_q0_1_166),
.o_LDPC_DEC_ERR_Q0_1_INTRO_167_err_intro_q0_1_167(o_LDPC_DEC_ERR_Q0_1_INTRO_167_err_intro_q0_1_167),
.o_LDPC_DEC_ERR_Q0_1_INTRO_168_err_intro_q0_1_168(o_LDPC_DEC_ERR_Q0_1_INTRO_168_err_intro_q0_1_168),
.o_LDPC_DEC_ERR_Q0_1_INTRO_169_err_intro_q0_1_169(o_LDPC_DEC_ERR_Q0_1_INTRO_169_err_intro_q0_1_169),
.o_LDPC_DEC_ERR_Q0_1_INTRO_170_err_intro_q0_1_170(o_LDPC_DEC_ERR_Q0_1_INTRO_170_err_intro_q0_1_170),
.o_LDPC_DEC_ERR_Q0_1_INTRO_171_err_intro_q0_1_171(o_LDPC_DEC_ERR_Q0_1_INTRO_171_err_intro_q0_1_171),
.o_LDPC_DEC_ERR_Q0_1_INTRO_172_err_intro_q0_1_172(o_LDPC_DEC_ERR_Q0_1_INTRO_172_err_intro_q0_1_172),
.o_LDPC_DEC_ERR_Q0_1_INTRO_173_err_intro_q0_1_173(o_LDPC_DEC_ERR_Q0_1_INTRO_173_err_intro_q0_1_173),
.o_LDPC_DEC_ERR_Q0_1_INTRO_174_err_intro_q0_1_174(o_LDPC_DEC_ERR_Q0_1_INTRO_174_err_intro_q0_1_174),
.o_LDPC_DEC_ERR_Q0_1_INTRO_175_err_intro_q0_1_175(o_LDPC_DEC_ERR_Q0_1_INTRO_175_err_intro_q0_1_175),
.o_LDPC_DEC_ERR_Q0_1_INTRO_176_err_intro_q0_1_176(o_LDPC_DEC_ERR_Q0_1_INTRO_176_err_intro_q0_1_176),
.o_LDPC_DEC_ERR_Q0_1_INTRO_177_err_intro_q0_1_177(o_LDPC_DEC_ERR_Q0_1_INTRO_177_err_intro_q0_1_177),
.o_LDPC_DEC_ERR_Q0_1_INTRO_178_err_intro_q0_1_178(o_LDPC_DEC_ERR_Q0_1_INTRO_178_err_intro_q0_1_178),
.o_LDPC_DEC_ERR_Q0_1_INTRO_179_err_intro_q0_1_179(o_LDPC_DEC_ERR_Q0_1_INTRO_179_err_intro_q0_1_179),
.o_LDPC_DEC_ERR_Q0_1_INTRO_180_err_intro_q0_1_180(o_LDPC_DEC_ERR_Q0_1_INTRO_180_err_intro_q0_1_180),
.o_LDPC_DEC_ERR_Q0_1_INTRO_181_err_intro_q0_1_181(o_LDPC_DEC_ERR_Q0_1_INTRO_181_err_intro_q0_1_181),
.o_LDPC_DEC_ERR_Q0_1_INTRO_182_err_intro_q0_1_182(o_LDPC_DEC_ERR_Q0_1_INTRO_182_err_intro_q0_1_182),
.o_LDPC_DEC_ERR_Q0_1_INTRO_183_err_intro_q0_1_183(o_LDPC_DEC_ERR_Q0_1_INTRO_183_err_intro_q0_1_183),
.o_LDPC_DEC_ERR_Q0_1_INTRO_184_err_intro_q0_1_184(o_LDPC_DEC_ERR_Q0_1_INTRO_184_err_intro_q0_1_184),
.o_LDPC_DEC_ERR_Q0_1_INTRO_185_err_intro_q0_1_185(o_LDPC_DEC_ERR_Q0_1_INTRO_185_err_intro_q0_1_185),
.o_LDPC_DEC_ERR_Q0_1_INTRO_186_err_intro_q0_1_186(o_LDPC_DEC_ERR_Q0_1_INTRO_186_err_intro_q0_1_186),
.o_LDPC_DEC_ERR_Q0_1_INTRO_187_err_intro_q0_1_187(o_LDPC_DEC_ERR_Q0_1_INTRO_187_err_intro_q0_1_187),
.o_LDPC_DEC_ERR_Q0_1_INTRO_188_err_intro_q0_1_188(o_LDPC_DEC_ERR_Q0_1_INTRO_188_err_intro_q0_1_188),
.o_LDPC_DEC_ERR_Q0_1_INTRO_189_err_intro_q0_1_189(o_LDPC_DEC_ERR_Q0_1_INTRO_189_err_intro_q0_1_189),
.o_LDPC_DEC_ERR_Q0_1_INTRO_190_err_intro_q0_1_190(o_LDPC_DEC_ERR_Q0_1_INTRO_190_err_intro_q0_1_190),
.o_LDPC_DEC_ERR_Q0_1_INTRO_191_err_intro_q0_1_191(o_LDPC_DEC_ERR_Q0_1_INTRO_191_err_intro_q0_1_191),
.o_LDPC_DEC_ERR_Q0_1_INTRO_192_err_intro_q0_1_192(o_LDPC_DEC_ERR_Q0_1_INTRO_192_err_intro_q0_1_192),
.o_LDPC_DEC_ERR_Q0_1_INTRO_193_err_intro_q0_1_193(o_LDPC_DEC_ERR_Q0_1_INTRO_193_err_intro_q0_1_193),
.o_LDPC_DEC_ERR_Q0_1_INTRO_194_err_intro_q0_1_194(o_LDPC_DEC_ERR_Q0_1_INTRO_194_err_intro_q0_1_194),
.o_LDPC_DEC_ERR_Q0_1_INTRO_195_err_intro_q0_1_195(o_LDPC_DEC_ERR_Q0_1_INTRO_195_err_intro_q0_1_195),
.o_LDPC_DEC_ERR_Q0_1_INTRO_196_err_intro_q0_1_196(o_LDPC_DEC_ERR_Q0_1_INTRO_196_err_intro_q0_1_196),
.o_LDPC_DEC_ERR_Q0_1_INTRO_197_err_intro_q0_1_197(o_LDPC_DEC_ERR_Q0_1_INTRO_197_err_intro_q0_1_197),
.o_LDPC_DEC_ERR_Q0_1_INTRO_198_err_intro_q0_1_198(o_LDPC_DEC_ERR_Q0_1_INTRO_198_err_intro_q0_1_198),
.o_LDPC_DEC_ERR_Q0_1_INTRO_199_err_intro_q0_1_199(o_LDPC_DEC_ERR_Q0_1_INTRO_199_err_intro_q0_1_199),
.o_LDPC_DEC_ERR_Q0_1_INTRO_200_err_intro_q0_1_200(o_LDPC_DEC_ERR_Q0_1_INTRO_200_err_intro_q0_1_200),
.o_LDPC_DEC_ERR_Q0_1_INTRO_201_err_intro_q0_1_201(o_LDPC_DEC_ERR_Q0_1_INTRO_201_err_intro_q0_1_201),
.o_LDPC_DEC_ERR_Q0_1_INTRO_202_err_intro_q0_1_202(o_LDPC_DEC_ERR_Q0_1_INTRO_202_err_intro_q0_1_202),
.o_LDPC_DEC_ERR_Q0_1_INTRO_203_err_intro_q0_1_203(o_LDPC_DEC_ERR_Q0_1_INTRO_203_err_intro_q0_1_203),
.o_LDPC_DEC_ERR_Q0_1_INTRO_204_err_intro_q0_1_204(o_LDPC_DEC_ERR_Q0_1_INTRO_204_err_intro_q0_1_204),
.o_LDPC_DEC_ERR_Q0_1_INTRO_205_err_intro_q0_1_205(o_LDPC_DEC_ERR_Q0_1_INTRO_205_err_intro_q0_1_205),
.o_LDPC_DEC_ERR_Q0_1_INTRO_206_err_intro_q0_1_206(o_LDPC_DEC_ERR_Q0_1_INTRO_206_err_intro_q0_1_206),
.o_LDPC_DEC_ERR_Q0_1_INTRO_207_err_intro_q0_1_207(o_LDPC_DEC_ERR_Q0_1_INTRO_207_err_intro_q0_1_207),
.o_LDPC_DEC_CODEWRD_IN_q0_0_0_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_0_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_1_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_1_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_2_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_2_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_3_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_3_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_4_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_4_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_5_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_5_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_6_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_6_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_7_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_7_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_8_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_8_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_9_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_9_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_10_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_10_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_11_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_11_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_12_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_12_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_13_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_13_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_14_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_14_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_15_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_15_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_16_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_16_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_17_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_17_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_18_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_18_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_19_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_19_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_20_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_20_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_21_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_21_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_22_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_22_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_23_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_23_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_24_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_24_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_25_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_25_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_26_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_26_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_27_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_27_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_28_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_28_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_29_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_29_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_30_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_30_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_31_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_31_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_32_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_32_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_33_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_33_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_34_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_34_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_35_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_35_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_36_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_36_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_37_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_37_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_38_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_38_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_39_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_39_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_40_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_40_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_41_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_41_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_42_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_42_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_43_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_43_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_44_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_44_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_45_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_45_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_46_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_46_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_47_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_47_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_48_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_48_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_49_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_49_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_50_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_50_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_51_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_51_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_52_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_52_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_53_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_53_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_54_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_54_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_55_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_55_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_56_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_56_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_57_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_57_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_58_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_58_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_59_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_59_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_60_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_60_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_61_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_61_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_62_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_62_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_63_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_63_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_64_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_64_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_65_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_65_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_66_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_66_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_67_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_67_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_68_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_68_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_69_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_69_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_70_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_70_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_71_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_71_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_72_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_72_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_73_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_73_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_74_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_74_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_75_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_75_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_76_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_76_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_77_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_77_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_78_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_78_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_79_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_79_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_80_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_80_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_81_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_81_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_82_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_82_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_83_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_83_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_84_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_84_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_85_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_85_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_86_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_86_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_87_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_87_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_88_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_88_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_89_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_89_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_90_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_90_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_91_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_91_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_92_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_92_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_93_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_93_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_94_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_94_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_95_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_95_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_96_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_96_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_97_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_97_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_98_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_98_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_99_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_99_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_100_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_100_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_101_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_101_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_102_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_102_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_103_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_103_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_104_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_104_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_105_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_105_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_106_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_106_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_107_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_107_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_108_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_108_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_109_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_109_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_110_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_110_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_111_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_111_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_112_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_112_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_113_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_113_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_114_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_114_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_115_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_115_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_116_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_116_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_117_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_117_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_118_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_118_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_119_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_119_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_120_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_120_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_121_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_121_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_122_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_122_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_123_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_123_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_124_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_124_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_125_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_125_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_126_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_126_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_127_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_127_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_128_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_128_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_129_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_129_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_130_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_130_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_131_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_131_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_132_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_132_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_133_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_133_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_134_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_134_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_135_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_135_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_136_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_136_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_137_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_137_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_138_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_138_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_139_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_139_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_140_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_140_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_141_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_141_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_142_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_142_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_143_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_143_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_144_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_144_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_145_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_145_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_146_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_146_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_147_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_147_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_148_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_148_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_149_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_149_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_150_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_150_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_151_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_151_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_152_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_152_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_153_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_153_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_154_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_154_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_155_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_155_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_156_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_156_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_157_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_157_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_158_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_158_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_159_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_159_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_160_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_160_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_161_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_161_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_162_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_162_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_163_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_163_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_164_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_164_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_165_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_165_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_166_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_166_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_167_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_167_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_168_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_168_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_169_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_169_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_170_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_170_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_171_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_171_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_172_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_172_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_173_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_173_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_174_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_174_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_175_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_175_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_176_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_176_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_177_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_177_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_178_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_178_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_179_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_179_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_180_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_180_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_181_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_181_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_182_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_182_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_183_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_183_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_184_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_184_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_185_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_185_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_186_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_186_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_187_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_187_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_188_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_188_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_189_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_189_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_190_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_190_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_191_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_191_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_192_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_192_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_193_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_193_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_194_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_194_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_195_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_195_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_196_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_196_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_197_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_197_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_198_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_198_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_199_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_199_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_200_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_200_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_201_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_201_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_202_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_202_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_203_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_203_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_204_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_204_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_205_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_205_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_206_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_206_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_0_207_cword_q0_0(o_LDPC_DEC_CODEWRD_IN_q0_0_207_cword_q0_0),
.o_LDPC_DEC_CODEWRD_IN_q0_1_0_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_0_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_1_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_1_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_2_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_2_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_3_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_3_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_4_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_4_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_5_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_5_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_6_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_6_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_7_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_7_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_8_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_8_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_9_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_9_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_10_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_10_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_11_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_11_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_12_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_12_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_13_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_13_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_14_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_14_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_15_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_15_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_16_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_16_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_17_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_17_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_18_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_18_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_19_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_19_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_20_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_20_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_21_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_21_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_22_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_22_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_23_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_23_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_24_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_24_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_25_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_25_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_26_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_26_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_27_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_27_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_28_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_28_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_29_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_29_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_30_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_30_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_31_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_31_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_32_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_32_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_33_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_33_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_34_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_34_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_35_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_35_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_36_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_36_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_37_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_37_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_38_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_38_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_39_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_39_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_40_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_40_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_41_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_41_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_42_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_42_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_43_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_43_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_44_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_44_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_45_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_45_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_46_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_46_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_47_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_47_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_48_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_48_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_49_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_49_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_50_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_50_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_51_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_51_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_52_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_52_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_53_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_53_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_54_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_54_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_55_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_55_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_56_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_56_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_57_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_57_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_58_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_58_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_59_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_59_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_60_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_60_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_61_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_61_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_62_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_62_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_63_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_63_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_64_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_64_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_65_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_65_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_66_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_66_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_67_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_67_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_68_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_68_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_69_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_69_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_70_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_70_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_71_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_71_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_72_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_72_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_73_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_73_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_74_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_74_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_75_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_75_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_76_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_76_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_77_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_77_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_78_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_78_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_79_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_79_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_80_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_80_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_81_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_81_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_82_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_82_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_83_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_83_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_84_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_84_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_85_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_85_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_86_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_86_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_87_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_87_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_88_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_88_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_89_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_89_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_90_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_90_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_91_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_91_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_92_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_92_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_93_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_93_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_94_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_94_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_95_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_95_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_96_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_96_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_97_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_97_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_98_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_98_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_99_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_99_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_100_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_100_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_101_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_101_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_102_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_102_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_103_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_103_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_104_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_104_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_105_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_105_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_106_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_106_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_107_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_107_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_108_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_108_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_109_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_109_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_110_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_110_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_111_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_111_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_112_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_112_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_113_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_113_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_114_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_114_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_115_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_115_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_116_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_116_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_117_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_117_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_118_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_118_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_119_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_119_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_120_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_120_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_121_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_121_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_122_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_122_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_123_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_123_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_124_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_124_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_125_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_125_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_126_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_126_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_127_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_127_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_128_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_128_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_129_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_129_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_130_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_130_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_131_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_131_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_132_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_132_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_133_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_133_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_134_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_134_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_135_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_135_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_136_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_136_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_137_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_137_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_138_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_138_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_139_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_139_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_140_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_140_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_141_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_141_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_142_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_142_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_143_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_143_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_144_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_144_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_145_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_145_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_146_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_146_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_147_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_147_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_148_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_148_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_149_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_149_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_150_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_150_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_151_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_151_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_152_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_152_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_153_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_153_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_154_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_154_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_155_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_155_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_156_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_156_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_157_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_157_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_158_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_158_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_159_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_159_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_160_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_160_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_161_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_161_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_162_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_162_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_163_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_163_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_164_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_164_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_165_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_165_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_166_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_166_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_167_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_167_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_168_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_168_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_169_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_169_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_170_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_170_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_171_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_171_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_172_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_172_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_173_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_173_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_174_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_174_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_175_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_175_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_176_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_176_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_177_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_177_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_178_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_178_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_179_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_179_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_180_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_180_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_181_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_181_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_182_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_182_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_183_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_183_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_184_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_184_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_185_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_185_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_186_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_186_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_187_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_187_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_188_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_188_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_189_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_189_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_190_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_190_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_191_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_191_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_192_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_192_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_193_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_193_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_194_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_194_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_195_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_195_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_196_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_196_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_197_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_197_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_198_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_198_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_199_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_199_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_200_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_200_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_201_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_201_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_202_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_202_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_203_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_203_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_204_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_204_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_205_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_205_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_206_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_206_cword_q0_1),
.o_LDPC_DEC_CODEWRD_IN_q0_1_207_cword_q0_1(o_LDPC_DEC_CODEWRD_IN_q0_1_207_cword_q0_1),
.i_LDPC_DEC_err_intro_decoder_err_intro_decoder_bit(i_LDPC_DEC_err_intro_decoder_err_intro_decoder_bit),
.o_LDPC_DEC_EXPSYND_0_exp_syn(o_LDPC_DEC_EXPSYND_0_exp_syn),
.o_LDPC_DEC_EXPSYND_1_exp_syn(o_LDPC_DEC_EXPSYND_1_exp_syn),
.o_LDPC_DEC_EXPSYND_2_exp_syn(o_LDPC_DEC_EXPSYND_2_exp_syn),
.o_LDPC_DEC_EXPSYND_3_exp_syn(o_LDPC_DEC_EXPSYND_3_exp_syn),
.o_LDPC_DEC_EXPSYND_4_exp_syn(o_LDPC_DEC_EXPSYND_4_exp_syn),
.o_LDPC_DEC_EXPSYND_5_exp_syn(o_LDPC_DEC_EXPSYND_5_exp_syn),
.o_LDPC_DEC_EXPSYND_6_exp_syn(o_LDPC_DEC_EXPSYND_6_exp_syn),
.o_LDPC_DEC_EXPSYND_7_exp_syn(o_LDPC_DEC_EXPSYND_7_exp_syn),
.o_LDPC_DEC_EXPSYND_8_exp_syn(o_LDPC_DEC_EXPSYND_8_exp_syn),
.o_LDPC_DEC_EXPSYND_9_exp_syn(o_LDPC_DEC_EXPSYND_9_exp_syn),
.o_LDPC_DEC_EXPSYND_10_exp_syn(o_LDPC_DEC_EXPSYND_10_exp_syn),
.o_LDPC_DEC_EXPSYND_11_exp_syn(o_LDPC_DEC_EXPSYND_11_exp_syn),
.o_LDPC_DEC_EXPSYND_12_exp_syn(o_LDPC_DEC_EXPSYND_12_exp_syn),
.o_LDPC_DEC_EXPSYND_13_exp_syn(o_LDPC_DEC_EXPSYND_13_exp_syn),
.o_LDPC_DEC_EXPSYND_14_exp_syn(o_LDPC_DEC_EXPSYND_14_exp_syn),
.o_LDPC_DEC_EXPSYND_15_exp_syn(o_LDPC_DEC_EXPSYND_15_exp_syn),
.o_LDPC_DEC_EXPSYND_16_exp_syn(o_LDPC_DEC_EXPSYND_16_exp_syn),
.o_LDPC_DEC_EXPSYND_17_exp_syn(o_LDPC_DEC_EXPSYND_17_exp_syn),
.o_LDPC_DEC_EXPSYND_18_exp_syn(o_LDPC_DEC_EXPSYND_18_exp_syn),
.o_LDPC_DEC_EXPSYND_19_exp_syn(o_LDPC_DEC_EXPSYND_19_exp_syn),
.o_LDPC_DEC_EXPSYND_20_exp_syn(o_LDPC_DEC_EXPSYND_20_exp_syn),
.o_LDPC_DEC_EXPSYND_21_exp_syn(o_LDPC_DEC_EXPSYND_21_exp_syn),
.o_LDPC_DEC_EXPSYND_22_exp_syn(o_LDPC_DEC_EXPSYND_22_exp_syn),
.o_LDPC_DEC_EXPSYND_23_exp_syn(o_LDPC_DEC_EXPSYND_23_exp_syn),
.o_LDPC_DEC_EXPSYND_24_exp_syn(o_LDPC_DEC_EXPSYND_24_exp_syn),
.o_LDPC_DEC_EXPSYND_25_exp_syn(o_LDPC_DEC_EXPSYND_25_exp_syn),
.o_LDPC_DEC_EXPSYND_26_exp_syn(o_LDPC_DEC_EXPSYND_26_exp_syn),
.o_LDPC_DEC_EXPSYND_27_exp_syn(o_LDPC_DEC_EXPSYND_27_exp_syn),
.o_LDPC_DEC_EXPSYND_28_exp_syn(o_LDPC_DEC_EXPSYND_28_exp_syn),
.o_LDPC_DEC_EXPSYND_29_exp_syn(o_LDPC_DEC_EXPSYND_29_exp_syn),
.o_LDPC_DEC_EXPSYND_30_exp_syn(o_LDPC_DEC_EXPSYND_30_exp_syn),
.o_LDPC_DEC_EXPSYND_31_exp_syn(o_LDPC_DEC_EXPSYND_31_exp_syn),
.o_LDPC_DEC_EXPSYND_32_exp_syn(o_LDPC_DEC_EXPSYND_32_exp_syn),
.o_LDPC_DEC_EXPSYND_33_exp_syn(o_LDPC_DEC_EXPSYND_33_exp_syn),
.o_LDPC_DEC_EXPSYND_34_exp_syn(o_LDPC_DEC_EXPSYND_34_exp_syn),
.o_LDPC_DEC_EXPSYND_35_exp_syn(o_LDPC_DEC_EXPSYND_35_exp_syn),
.o_LDPC_DEC_EXPSYND_36_exp_syn(o_LDPC_DEC_EXPSYND_36_exp_syn),
.o_LDPC_DEC_EXPSYND_37_exp_syn(o_LDPC_DEC_EXPSYND_37_exp_syn),
.o_LDPC_DEC_EXPSYND_38_exp_syn(o_LDPC_DEC_EXPSYND_38_exp_syn),
.o_LDPC_DEC_EXPSYND_39_exp_syn(o_LDPC_DEC_EXPSYND_39_exp_syn),
.o_LDPC_DEC_EXPSYND_40_exp_syn(o_LDPC_DEC_EXPSYND_40_exp_syn),
.o_LDPC_DEC_EXPSYND_41_exp_syn(o_LDPC_DEC_EXPSYND_41_exp_syn),
.o_LDPC_DEC_EXPSYND_42_exp_syn(o_LDPC_DEC_EXPSYND_42_exp_syn),
.o_LDPC_DEC_EXPSYND_43_exp_syn(o_LDPC_DEC_EXPSYND_43_exp_syn),
.o_LDPC_DEC_EXPSYND_44_exp_syn(o_LDPC_DEC_EXPSYND_44_exp_syn),
.o_LDPC_DEC_EXPSYND_45_exp_syn(o_LDPC_DEC_EXPSYND_45_exp_syn),
.o_LDPC_DEC_EXPSYND_46_exp_syn(o_LDPC_DEC_EXPSYND_46_exp_syn),
.o_LDPC_DEC_EXPSYND_47_exp_syn(o_LDPC_DEC_EXPSYND_47_exp_syn),
.o_LDPC_DEC_EXPSYND_48_exp_syn(o_LDPC_DEC_EXPSYND_48_exp_syn),
.o_LDPC_DEC_EXPSYND_49_exp_syn(o_LDPC_DEC_EXPSYND_49_exp_syn),
.o_LDPC_DEC_EXPSYND_50_exp_syn(o_LDPC_DEC_EXPSYND_50_exp_syn),
.o_LDPC_DEC_EXPSYND_51_exp_syn(o_LDPC_DEC_EXPSYND_51_exp_syn),
.o_LDPC_DEC_EXPSYND_52_exp_syn(o_LDPC_DEC_EXPSYND_52_exp_syn),
.o_LDPC_DEC_EXPSYND_53_exp_syn(o_LDPC_DEC_EXPSYND_53_exp_syn),
.o_LDPC_DEC_EXPSYND_54_exp_syn(o_LDPC_DEC_EXPSYND_54_exp_syn),
.o_LDPC_DEC_EXPSYND_55_exp_syn(o_LDPC_DEC_EXPSYND_55_exp_syn),
.o_LDPC_DEC_EXPSYND_56_exp_syn(o_LDPC_DEC_EXPSYND_56_exp_syn),
.o_LDPC_DEC_EXPSYND_57_exp_syn(o_LDPC_DEC_EXPSYND_57_exp_syn),
.o_LDPC_DEC_EXPSYND_58_exp_syn(o_LDPC_DEC_EXPSYND_58_exp_syn),
.o_LDPC_DEC_EXPSYND_59_exp_syn(o_LDPC_DEC_EXPSYND_59_exp_syn),
.o_LDPC_DEC_EXPSYND_60_exp_syn(o_LDPC_DEC_EXPSYND_60_exp_syn),
.o_LDPC_DEC_EXPSYND_61_exp_syn(o_LDPC_DEC_EXPSYND_61_exp_syn),
.o_LDPC_DEC_EXPSYND_62_exp_syn(o_LDPC_DEC_EXPSYND_62_exp_syn),
.o_LDPC_DEC_EXPSYND_63_exp_syn(o_LDPC_DEC_EXPSYND_63_exp_syn),
.o_LDPC_DEC_EXPSYND_64_exp_syn(o_LDPC_DEC_EXPSYND_64_exp_syn),
.o_LDPC_DEC_EXPSYND_65_exp_syn(o_LDPC_DEC_EXPSYND_65_exp_syn),
.o_LDPC_DEC_EXPSYND_66_exp_syn(o_LDPC_DEC_EXPSYND_66_exp_syn),
.o_LDPC_DEC_EXPSYND_67_exp_syn(o_LDPC_DEC_EXPSYND_67_exp_syn),
.o_LDPC_DEC_EXPSYND_68_exp_syn(o_LDPC_DEC_EXPSYND_68_exp_syn),
.o_LDPC_DEC_EXPSYND_69_exp_syn(o_LDPC_DEC_EXPSYND_69_exp_syn),
.o_LDPC_DEC_EXPSYND_70_exp_syn(o_LDPC_DEC_EXPSYND_70_exp_syn),
.o_LDPC_DEC_EXPSYND_71_exp_syn(o_LDPC_DEC_EXPSYND_71_exp_syn),
.o_LDPC_DEC_EXPSYND_72_exp_syn(o_LDPC_DEC_EXPSYND_72_exp_syn),
.o_LDPC_DEC_EXPSYND_73_exp_syn(o_LDPC_DEC_EXPSYND_73_exp_syn),
.o_LDPC_DEC_EXPSYND_74_exp_syn(o_LDPC_DEC_EXPSYND_74_exp_syn),
.o_LDPC_DEC_EXPSYND_75_exp_syn(o_LDPC_DEC_EXPSYND_75_exp_syn),
.o_LDPC_DEC_EXPSYND_76_exp_syn(o_LDPC_DEC_EXPSYND_76_exp_syn),
.o_LDPC_DEC_EXPSYND_77_exp_syn(o_LDPC_DEC_EXPSYND_77_exp_syn),
.o_LDPC_DEC_EXPSYND_78_exp_syn(o_LDPC_DEC_EXPSYND_78_exp_syn),
.o_LDPC_DEC_EXPSYND_79_exp_syn(o_LDPC_DEC_EXPSYND_79_exp_syn),
.o_LDPC_DEC_EXPSYND_80_exp_syn(o_LDPC_DEC_EXPSYND_80_exp_syn),
.o_LDPC_DEC_EXPSYND_81_exp_syn(o_LDPC_DEC_EXPSYND_81_exp_syn),
.o_LDPC_DEC_EXPSYND_82_exp_syn(o_LDPC_DEC_EXPSYND_82_exp_syn),
.o_LDPC_DEC_EXPSYND_83_exp_syn(o_LDPC_DEC_EXPSYND_83_exp_syn),
.o_LDPC_DEC_EXPSYND_84_exp_syn(o_LDPC_DEC_EXPSYND_84_exp_syn),
.o_LDPC_DEC_EXPSYND_85_exp_syn(o_LDPC_DEC_EXPSYND_85_exp_syn),
.o_LDPC_DEC_EXPSYND_86_exp_syn(o_LDPC_DEC_EXPSYND_86_exp_syn),
.o_LDPC_DEC_EXPSYND_87_exp_syn(o_LDPC_DEC_EXPSYND_87_exp_syn),
.o_LDPC_DEC_EXPSYND_88_exp_syn(o_LDPC_DEC_EXPSYND_88_exp_syn),
.o_LDPC_DEC_EXPSYND_89_exp_syn(o_LDPC_DEC_EXPSYND_89_exp_syn),
.o_LDPC_DEC_EXPSYND_90_exp_syn(o_LDPC_DEC_EXPSYND_90_exp_syn),
.o_LDPC_DEC_EXPSYND_91_exp_syn(o_LDPC_DEC_EXPSYND_91_exp_syn),
.o_LDPC_DEC_EXPSYND_92_exp_syn(o_LDPC_DEC_EXPSYND_92_exp_syn),
.o_LDPC_DEC_EXPSYND_93_exp_syn(o_LDPC_DEC_EXPSYND_93_exp_syn),
.o_LDPC_DEC_EXPSYND_94_exp_syn(o_LDPC_DEC_EXPSYND_94_exp_syn),
.o_LDPC_DEC_EXPSYND_95_exp_syn(o_LDPC_DEC_EXPSYND_95_exp_syn),
.o_LDPC_DEC_EXPSYND_96_exp_syn(o_LDPC_DEC_EXPSYND_96_exp_syn),
.o_LDPC_DEC_EXPSYND_97_exp_syn(o_LDPC_DEC_EXPSYND_97_exp_syn),
.o_LDPC_DEC_EXPSYND_98_exp_syn(o_LDPC_DEC_EXPSYND_98_exp_syn),
.o_LDPC_DEC_EXPSYND_99_exp_syn(o_LDPC_DEC_EXPSYND_99_exp_syn),
.o_LDPC_DEC_EXPSYND_100_exp_syn(o_LDPC_DEC_EXPSYND_100_exp_syn),
.o_LDPC_DEC_EXPSYND_101_exp_syn(o_LDPC_DEC_EXPSYND_101_exp_syn),
.o_LDPC_DEC_EXPSYND_102_exp_syn(o_LDPC_DEC_EXPSYND_102_exp_syn),
.o_LDPC_DEC_EXPSYND_103_exp_syn(o_LDPC_DEC_EXPSYND_103_exp_syn),
.o_LDPC_DEC_EXPSYND_104_exp_syn(o_LDPC_DEC_EXPSYND_104_exp_syn),
.o_LDPC_DEC_EXPSYND_105_exp_syn(o_LDPC_DEC_EXPSYND_105_exp_syn),
.o_LDPC_DEC_EXPSYND_106_exp_syn(o_LDPC_DEC_EXPSYND_106_exp_syn),
.o_LDPC_DEC_EXPSYND_107_exp_syn(o_LDPC_DEC_EXPSYND_107_exp_syn),
.o_LDPC_DEC_EXPSYND_108_exp_syn(o_LDPC_DEC_EXPSYND_108_exp_syn),
.o_LDPC_DEC_EXPSYND_109_exp_syn(o_LDPC_DEC_EXPSYND_109_exp_syn),
.o_LDPC_DEC_EXPSYND_110_exp_syn(o_LDPC_DEC_EXPSYND_110_exp_syn),
.o_LDPC_DEC_EXPSYND_111_exp_syn(o_LDPC_DEC_EXPSYND_111_exp_syn),
.o_LDPC_DEC_EXPSYND_112_exp_syn(o_LDPC_DEC_EXPSYND_112_exp_syn),
.o_LDPC_DEC_EXPSYND_113_exp_syn(o_LDPC_DEC_EXPSYND_113_exp_syn),
.o_LDPC_DEC_EXPSYND_114_exp_syn(o_LDPC_DEC_EXPSYND_114_exp_syn),
.o_LDPC_DEC_EXPSYND_115_exp_syn(o_LDPC_DEC_EXPSYND_115_exp_syn),
.o_LDPC_DEC_EXPSYND_116_exp_syn(o_LDPC_DEC_EXPSYND_116_exp_syn),
.o_LDPC_DEC_EXPSYND_117_exp_syn(o_LDPC_DEC_EXPSYND_117_exp_syn),
.o_LDPC_DEC_EXPSYND_118_exp_syn(o_LDPC_DEC_EXPSYND_118_exp_syn),
.o_LDPC_DEC_EXPSYND_119_exp_syn(o_LDPC_DEC_EXPSYND_119_exp_syn),
.o_LDPC_DEC_EXPSYND_120_exp_syn(o_LDPC_DEC_EXPSYND_120_exp_syn),
.o_LDPC_DEC_EXPSYND_121_exp_syn(o_LDPC_DEC_EXPSYND_121_exp_syn),
.o_LDPC_DEC_EXPSYND_122_exp_syn(o_LDPC_DEC_EXPSYND_122_exp_syn),
.o_LDPC_DEC_EXPSYND_123_exp_syn(o_LDPC_DEC_EXPSYND_123_exp_syn),
.o_LDPC_DEC_EXPSYND_124_exp_syn(o_LDPC_DEC_EXPSYND_124_exp_syn),
.o_LDPC_DEC_EXPSYND_125_exp_syn(o_LDPC_DEC_EXPSYND_125_exp_syn),
.o_LDPC_DEC_EXPSYND_126_exp_syn(o_LDPC_DEC_EXPSYND_126_exp_syn),
.o_LDPC_DEC_EXPSYND_127_exp_syn(o_LDPC_DEC_EXPSYND_127_exp_syn),
.o_LDPC_DEC_EXPSYND_128_exp_syn(o_LDPC_DEC_EXPSYND_128_exp_syn),
.o_LDPC_DEC_EXPSYND_129_exp_syn(o_LDPC_DEC_EXPSYND_129_exp_syn),
.o_LDPC_DEC_EXPSYND_130_exp_syn(o_LDPC_DEC_EXPSYND_130_exp_syn),
.o_LDPC_DEC_EXPSYND_131_exp_syn(o_LDPC_DEC_EXPSYND_131_exp_syn),
.o_LDPC_DEC_EXPSYND_132_exp_syn(o_LDPC_DEC_EXPSYND_132_exp_syn),
.o_LDPC_DEC_EXPSYND_133_exp_syn(o_LDPC_DEC_EXPSYND_133_exp_syn),
.o_LDPC_DEC_EXPSYND_134_exp_syn(o_LDPC_DEC_EXPSYND_134_exp_syn),
.o_LDPC_DEC_EXPSYND_135_exp_syn(o_LDPC_DEC_EXPSYND_135_exp_syn),
.o_LDPC_DEC_EXPSYND_136_exp_syn(o_LDPC_DEC_EXPSYND_136_exp_syn),
.o_LDPC_DEC_EXPSYND_137_exp_syn(o_LDPC_DEC_EXPSYND_137_exp_syn),
.o_LDPC_DEC_EXPSYND_138_exp_syn(o_LDPC_DEC_EXPSYND_138_exp_syn),
.o_LDPC_DEC_EXPSYND_139_exp_syn(o_LDPC_DEC_EXPSYND_139_exp_syn),
.o_LDPC_DEC_EXPSYND_140_exp_syn(o_LDPC_DEC_EXPSYND_140_exp_syn),
.o_LDPC_DEC_EXPSYND_141_exp_syn(o_LDPC_DEC_EXPSYND_141_exp_syn),
.o_LDPC_DEC_EXPSYND_142_exp_syn(o_LDPC_DEC_EXPSYND_142_exp_syn),
.o_LDPC_DEC_EXPSYND_143_exp_syn(o_LDPC_DEC_EXPSYND_143_exp_syn),
.o_LDPC_DEC_EXPSYND_144_exp_syn(o_LDPC_DEC_EXPSYND_144_exp_syn),
.o_LDPC_DEC_EXPSYND_145_exp_syn(o_LDPC_DEC_EXPSYND_145_exp_syn),
.o_LDPC_DEC_EXPSYND_146_exp_syn(o_LDPC_DEC_EXPSYND_146_exp_syn),
.o_LDPC_DEC_EXPSYND_147_exp_syn(o_LDPC_DEC_EXPSYND_147_exp_syn),
.o_LDPC_DEC_EXPSYND_148_exp_syn(o_LDPC_DEC_EXPSYND_148_exp_syn),
.o_LDPC_DEC_EXPSYND_149_exp_syn(o_LDPC_DEC_EXPSYND_149_exp_syn),
.o_LDPC_DEC_EXPSYND_150_exp_syn(o_LDPC_DEC_EXPSYND_150_exp_syn),
.o_LDPC_DEC_EXPSYND_151_exp_syn(o_LDPC_DEC_EXPSYND_151_exp_syn),
.o_LDPC_DEC_EXPSYND_152_exp_syn(o_LDPC_DEC_EXPSYND_152_exp_syn),
.o_LDPC_DEC_EXPSYND_153_exp_syn(o_LDPC_DEC_EXPSYND_153_exp_syn),
.o_LDPC_DEC_EXPSYND_154_exp_syn(o_LDPC_DEC_EXPSYND_154_exp_syn),
.o_LDPC_DEC_EXPSYND_155_exp_syn(o_LDPC_DEC_EXPSYND_155_exp_syn),
.o_LDPC_DEC_EXPSYND_156_exp_syn(o_LDPC_DEC_EXPSYND_156_exp_syn),
.o_LDPC_DEC_EXPSYND_157_exp_syn(o_LDPC_DEC_EXPSYND_157_exp_syn),
.o_LDPC_DEC_EXPSYND_158_exp_syn(o_LDPC_DEC_EXPSYND_158_exp_syn),
.o_LDPC_DEC_EXPSYND_159_exp_syn(o_LDPC_DEC_EXPSYND_159_exp_syn),
.o_LDPC_DEC_EXPSYND_160_exp_syn(o_LDPC_DEC_EXPSYND_160_exp_syn),
.o_LDPC_DEC_EXPSYND_161_exp_syn(o_LDPC_DEC_EXPSYND_161_exp_syn),
.o_LDPC_DEC_EXPSYND_162_exp_syn(o_LDPC_DEC_EXPSYND_162_exp_syn),
.o_LDPC_DEC_EXPSYND_163_exp_syn(o_LDPC_DEC_EXPSYND_163_exp_syn),
.o_LDPC_DEC_EXPSYND_164_exp_syn(o_LDPC_DEC_EXPSYND_164_exp_syn),
.o_LDPC_DEC_EXPSYND_165_exp_syn(o_LDPC_DEC_EXPSYND_165_exp_syn),
.o_LDPC_DEC_EXPSYND_166_exp_syn(o_LDPC_DEC_EXPSYND_166_exp_syn),
.o_LDPC_DEC_EXPSYND_167_exp_syn(o_LDPC_DEC_EXPSYND_167_exp_syn),
.o_LDPC_DEC_PROBABILITY_perc_probability(o_LDPC_DEC_PROBABILITY_perc_probability),
.o_LDPC_DEC_HAMDIST_LOOP_MAX_HamDist_loop_max(o_LDPC_DEC_HAMDIST_LOOP_MAX_HamDist_loop_max),
.o_LDPC_DEC_HAMDIST_LOOP_PERCENTAGE_HamDist_loop_percentage(o_LDPC_DEC_HAMDIST_LOOP_PERCENTAGE_HamDist_loop_percentage),
.o_LDPC_DEC_HAMDIST_IIR1_HamDist_iir1(o_LDPC_DEC_HAMDIST_IIR1_HamDist_iir1),
.o_LDPC_DEC_HAMDIST_IIR2_NOT_USED_HamDist_iir2(o_LDPC_DEC_HAMDIST_IIR2_NOT_USED_HamDist_iir2),
.o_LDPC_DEC_HAMDIST_IIR3_NOT_USED_HamDist_iir3(o_LDPC_DEC_HAMDIST_IIR3_NOT_USED_HamDist_iir3),
.i_LDPC_DEC_SYN_VALID_CWORD_DEC_final_syn_valid_cword_dec(i_LDPC_DEC_SYN_VALID_CWORD_DEC_final_syn_valid_cword_dec),
.o_LDPC_DEC_START_DEC_start_dec(o_LDPC_DEC_START_DEC_start_dec),
.i_LDPC_DEC_CONVERGED_LOOPS_ENDED_converged_loops_ended(i_LDPC_DEC_CONVERGED_LOOPS_ENDED_converged_loops_ended),
.i_LDPC_DEC_CONVERGED_PASS_FAIL_converged_pass_fail(i_LDPC_DEC_CONVERGED_PASS_FAIL_converged_pass_fail),
.i_LDPC_DEC_CODEWRD_OUT_BIT_0_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_0_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_1_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_1_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_2_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_2_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_3_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_3_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_4_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_4_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_5_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_5_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_6_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_6_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_7_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_7_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_8_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_8_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_9_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_9_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_10_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_10_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_11_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_11_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_12_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_12_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_13_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_13_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_14_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_14_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_15_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_15_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_16_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_16_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_17_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_17_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_18_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_18_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_19_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_19_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_20_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_20_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_21_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_21_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_22_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_22_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_23_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_23_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_24_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_24_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_25_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_25_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_26_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_26_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_27_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_27_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_28_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_28_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_29_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_29_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_30_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_30_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_31_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_31_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_32_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_32_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_33_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_33_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_34_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_34_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_35_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_35_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_36_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_36_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_37_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_37_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_38_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_38_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_39_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_39_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_40_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_40_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_41_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_41_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_42_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_42_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_43_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_43_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_44_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_44_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_45_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_45_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_46_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_46_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_47_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_47_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_48_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_48_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_49_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_49_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_50_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_50_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_51_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_51_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_52_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_52_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_53_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_53_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_54_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_54_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_55_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_55_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_56_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_56_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_57_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_57_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_58_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_58_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_59_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_59_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_60_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_60_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_61_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_61_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_62_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_62_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_63_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_63_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_64_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_64_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_65_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_65_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_66_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_66_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_67_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_67_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_68_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_68_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_69_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_69_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_70_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_70_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_71_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_71_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_72_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_72_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_73_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_73_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_74_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_74_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_75_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_75_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_76_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_76_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_77_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_77_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_78_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_78_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_79_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_79_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_80_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_80_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_81_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_81_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_82_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_82_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_83_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_83_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_84_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_84_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_85_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_85_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_86_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_86_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_87_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_87_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_88_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_88_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_89_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_89_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_90_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_90_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_91_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_91_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_92_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_92_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_93_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_93_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_94_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_94_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_95_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_95_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_96_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_96_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_97_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_97_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_98_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_98_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_99_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_99_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_100_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_100_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_101_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_101_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_102_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_102_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_103_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_103_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_104_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_104_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_105_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_105_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_106_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_106_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_107_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_107_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_108_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_108_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_109_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_109_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_110_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_110_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_111_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_111_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_112_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_112_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_113_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_113_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_114_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_114_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_115_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_115_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_116_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_116_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_117_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_117_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_118_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_118_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_119_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_119_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_120_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_120_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_121_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_121_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_122_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_122_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_123_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_123_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_124_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_124_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_125_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_125_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_126_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_126_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_127_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_127_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_128_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_128_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_129_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_129_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_130_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_130_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_131_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_131_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_132_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_132_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_133_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_133_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_134_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_134_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_135_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_135_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_136_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_136_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_137_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_137_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_138_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_138_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_139_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_139_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_140_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_140_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_141_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_141_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_142_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_142_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_143_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_143_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_144_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_144_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_145_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_145_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_146_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_146_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_147_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_147_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_148_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_148_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_149_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_149_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_150_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_150_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_151_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_151_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_152_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_152_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_153_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_153_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_154_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_154_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_155_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_155_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_156_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_156_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_157_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_157_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_158_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_158_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_159_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_159_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_160_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_160_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_161_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_161_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_162_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_162_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_163_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_163_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_164_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_164_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_165_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_165_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_166_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_166_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_167_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_167_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_168_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_168_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_169_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_169_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_170_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_170_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_171_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_171_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_172_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_172_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_173_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_173_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_174_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_174_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_175_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_175_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_176_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_176_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_177_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_177_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_178_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_178_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_179_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_179_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_180_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_180_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_181_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_181_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_182_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_182_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_183_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_183_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_184_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_184_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_185_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_185_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_186_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_186_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_187_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_187_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_188_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_188_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_189_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_189_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_190_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_190_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_191_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_191_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_192_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_192_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_193_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_193_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_194_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_194_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_195_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_195_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_196_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_196_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_197_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_197_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_198_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_198_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_199_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_199_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_200_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_200_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_201_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_201_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_202_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_202_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_203_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_203_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_204_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_204_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_205_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_205_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_206_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_206_final_cword),
.i_LDPC_DEC_CODEWRD_OUT_BIT_207_final_cword(i_LDPC_DEC_CODEWRD_OUT_BIT_207_final_cword),
.o_LDPC_DEC_PASS_FAIL_pass_fail(o_LDPC_DEC_PASS_FAIL_pass_fail),
.i_LDPC_DEC_pass_fail_decoder_pass_fail_decoder_bit(i_LDPC_DEC_pass_fail_decoder_pass_fail_decoder_bit),
