              fgallag0x00005_0 = 
          (!fgallag_sel[4]) ? 
                       fgallag0x00004_0_q: 
                       fgallag0x00004_1_q;
              fgallag0x00005_1 = 
          (!fgallag_sel[4]) ? 
                       fgallag0x00004_2_q: 
                       fgallag0x00004_3_q;
              fgallag0x00005_2 = 
          (!fgallag_sel[4]) ? 
                       fgallag0x00004_4_q: 
                       fgallag0x00004_5_q;
              fgallag0x00005_3 = 
          (!fgallag_sel[4]) ? 
                       fgallag0x00004_6_q: 
                       fgallag0x00004_7_q;
              fgallag0x00005_4 = 
          (!fgallag_sel[4]) ? 
                       fgallag0x00004_8_q: 
                       fgallag0x00004_9_q;
              fgallag0x00005_5 = 
          (!fgallag_sel[4]) ? 
                       fgallag0x00004_10_q: 
                       fgallag0x00004_11_q;
              fgallag0x00005_6 = 
          (!fgallag_sel[4]) ? 
                       fgallag0x00004_12_q: 
                       fgallag0x00004_13_q;
              fgallag0x00005_7 = 
          (!fgallag_sel[4]) ? 
                       fgallag0x00004_14_q: 
                       fgallag0x00004_15_q;
              fgallag0x00005_8 = 
          (!fgallag_sel[4]) ? 
                       fgallag0x00004_16_q: 
                       fgallag0x00004_17_q;
               fgallag0x00005_9 =  fgallag0x00004_18_q ;
               fgallag0x00005_10 =  fgallag0x00004_20_q ;
              fgallag0x00005_11 = 
          (!fgallag_sel[4]) ? 
                       fgallag0x00004_22_q: 
                       fgallag0x00004_23_q;
