              flogtanh0x00005_0 = 
          (!flogtanh_sel[4]) ? 
                       flogtanh0x00004_0_q: 
                       flogtanh0x00004_1_q;
              flogtanh0x00005_1 = 
          (!flogtanh_sel[4]) ? 
                       flogtanh0x00004_2_q: 
                       flogtanh0x00004_3_q;
              flogtanh0x00005_2 = 
          (!flogtanh_sel[4]) ? 
                       flogtanh0x00004_4_q: 
                       flogtanh0x00004_5_q;
              flogtanh0x00005_3 = 
          (!flogtanh_sel[4]) ? 
                       flogtanh0x00004_6_q: 
                       flogtanh0x00004_7_q;
              flogtanh0x00005_4 = 
          (!flogtanh_sel[4]) ? 
                       flogtanh0x00004_8_q: 
                       flogtanh0x00004_9_q;
              flogtanh0x00005_5 = 
          (!flogtanh_sel[4]) ? 
                       flogtanh0x00004_10_q: 
                       flogtanh0x00004_11_q;
              flogtanh0x00005_6 = 
          (!flogtanh_sel[4]) ? 
                       flogtanh0x00004_12_q: 
                       flogtanh0x00004_13_q;
              flogtanh0x00005_7 = 
          (!flogtanh_sel[4]) ? 
                       flogtanh0x00004_14_q: 
                       flogtanh0x00004_15_q;
              flogtanh0x00005_8 = 
          (!flogtanh_sel[4]) ? 
                       flogtanh0x00004_16_q: 
                       flogtanh0x00004_17_q;
               flogtanh0x00005_9 =  flogtanh0x00004_18_q ;
               flogtanh0x00005_10 =  flogtanh0x00004_20_q ;
              flogtanh0x00005_11 = 
          (!flogtanh_sel[4]) ? 
                       flogtanh0x00004_22_q: 
                       flogtanh0x00004_23_q;
