              fgallag0x00001_0 = 
          (!fgallag_sel[0]) ? 
                       fgallag0x00000_0_q: 
                       fgallag0x00000_1_q;
              fgallag0x00001_1 = 
          (!fgallag_sel[0]) ? 
                       fgallag0x00000_2_q: 
                       fgallag0x00000_3_q;
              fgallag0x00001_2 = 
          (!fgallag_sel[0]) ? 
                       fgallag0x00000_4_q: 
                       fgallag0x00000_5_q;
              fgallag0x00001_3 = 
          (!fgallag_sel[0]) ? 
                       fgallag0x00000_6_q: 
                       fgallag0x00000_7_q;
              fgallag0x00001_4 = 
          (!fgallag_sel[0]) ? 
                       fgallag0x00000_8_q: 
                       fgallag0x00000_9_q;
              fgallag0x00001_5 = 
          (!fgallag_sel[0]) ? 
                       fgallag0x00000_10_q: 
                       fgallag0x00000_11_q;
              fgallag0x00001_6 = 
          (!fgallag_sel[0]) ? 
                       fgallag0x00000_12_q: 
                       fgallag0x00000_13_q;
              fgallag0x00001_7 = 
          (!fgallag_sel[0]) ? 
                       fgallag0x00000_14_q: 
                       fgallag0x00000_15_q;
              fgallag0x00001_8 = 
          (!fgallag_sel[0]) ? 
                       fgallag0x00000_16_q: 
                       fgallag0x00000_17_q;
              fgallag0x00001_9 = 
          (!fgallag_sel[0]) ? 
                       fgallag0x00000_18_q: 
                       fgallag0x00000_19_q;
              fgallag0x00001_10 = 
          (!fgallag_sel[0]) ? 
                       fgallag0x00000_20_q: 
                       fgallag0x00000_21_q;
              fgallag0x00001_11 = 
          (!fgallag_sel[0]) ? 
                       fgallag0x00000_22_q: 
                       fgallag0x00000_23_q;
              fgallag0x00001_12 = 
          (!fgallag_sel[0]) ? 
                       fgallag0x00000_24_q: 
                       fgallag0x00000_25_q;
              fgallag0x00001_13 = 
          (!fgallag_sel[0]) ? 
                       fgallag0x00000_26_q: 
                       fgallag0x00000_27_q;
              fgallag0x00001_14 = 
          (!fgallag_sel[0]) ? 
                       fgallag0x00000_28_q: 
                       fgallag0x00000_29_q;
              fgallag0x00001_15 = 
          (!fgallag_sel[0]) ? 
                       fgallag0x00000_30_q: 
                       fgallag0x00000_31_q;
              fgallag0x00001_16 = 
          (!fgallag_sel[0]) ? 
                       fgallag0x00000_32_q: 
                       fgallag0x00000_33_q;
              fgallag0x00001_17 = 
          (!fgallag_sel[0]) ? 
                       fgallag0x00000_34_q: 
                       fgallag0x00000_35_q;
              fgallag0x00001_18 = 
          (!fgallag_sel[0]) ? 
                       fgallag0x00000_36_q: 
                       fgallag0x00000_37_q;
              fgallag0x00001_19 = 
          (!fgallag_sel[0]) ? 
                       fgallag0x00000_38_q: 
                       fgallag0x00000_39_q;
              fgallag0x00001_20 = 
          (!fgallag_sel[0]) ? 
                       fgallag0x00000_40_q: 
                       fgallag0x00000_41_q;
              fgallag0x00001_21 = 
          (!fgallag_sel[0]) ? 
                       fgallag0x00000_42_q: 
                       fgallag0x00000_43_q;
              fgallag0x00001_22 = 
          (!fgallag_sel[0]) ? 
                       fgallag0x00000_44_q: 
                       fgallag0x00000_45_q;
              fgallag0x00001_23 = 
          (!fgallag_sel[0]) ? 
                       fgallag0x00000_46_q: 
                       fgallag0x00000_47_q;
              fgallag0x00001_24 = 
          (!fgallag_sel[0]) ? 
                       fgallag0x00000_48_q: 
                       fgallag0x00000_49_q;
              fgallag0x00001_25 = 
          (!fgallag_sel[0]) ? 
                       fgallag0x00000_50_q: 
                       fgallag0x00000_51_q;
              fgallag0x00001_26 = 
          (!fgallag_sel[0]) ? 
                       fgallag0x00000_52_q: 
                       fgallag0x00000_53_q;
              fgallag0x00001_27 = 
          (!fgallag_sel[0]) ? 
                       fgallag0x00000_54_q: 
                       fgallag0x00000_55_q;
              fgallag0x00001_28 = 
          (!fgallag_sel[0]) ? 
                       fgallag0x00000_56_q: 
                       fgallag0x00000_57_q;
              fgallag0x00001_29 = 
          (!fgallag_sel[0]) ? 
                       fgallag0x00000_58_q: 
                       fgallag0x00000_59_q;
              fgallag0x00001_30 = 
          (!fgallag_sel[0]) ? 
                       fgallag0x00000_60_q: 
                       fgallag0x00000_61_q;
               fgallag0x00001_31 =  fgallag0x00000_62_q ;
              fgallag0x00001_32 = 
          (!fgallag_sel[0]) ? 
                       fgallag0x00000_64_q: 
                       fgallag0x00000_65_q;
              fgallag0x00001_33 = 
          (!fgallag_sel[0]) ? 
                       fgallag0x00000_66_q: 
                       fgallag0x00000_67_q;
               fgallag0x00001_34 =  fgallag0x00000_68_q ;
              fgallag0x00001_35 = 
          (!fgallag_sel[0]) ? 
                       fgallag0x00000_70_q: 
                       fgallag0x00000_71_q;
               fgallag0x00001_36 =  fgallag0x00000_72_q ;
              fgallag0x00001_37 = 
          (!fgallag_sel[0]) ? 
                       fgallag0x00000_74_q: 
                       fgallag0x00000_75_q;
              fgallag0x00001_38 = 
          (!fgallag_sel[0]) ? 
                       fgallag0x00000_76_q: 
                       fgallag0x00000_77_q;
               fgallag0x00001_39 =  fgallag0x00000_78_q ;
              fgallag0x00001_40 = 
          (!fgallag_sel[0]) ? 
                       fgallag0x00000_80_q: 
                       fgallag0x00000_81_q;
              fgallag0x00001_41 = 
          (!fgallag_sel[0]) ? 
                       fgallag0x00000_82_q: 
                       fgallag0x00000_83_q;
              fgallag0x00001_42 = 
          (!fgallag_sel[0]) ? 
                       fgallag0x00000_84_q: 
                       fgallag0x00000_85_q;
               fgallag0x00001_43 =  fgallag0x00000_86_q ;
               fgallag0x00001_44 =  fgallag0x00000_88_q ;
               fgallag0x00001_45 =  fgallag0x00000_90_q ;
               fgallag0x00001_46 =  fgallag0x00000_92_q ;
               fgallag0x00001_47 =  fgallag0x00000_94_q ;
               fgallag0x00001_48 =  fgallag0x00000_96_q ;
               fgallag0x00001_49 =  fgallag0x00000_98_q ;
               fgallag0x00001_50 =  fgallag0x00000_100_q ;
              fgallag0x00001_51 = 
          (!fgallag_sel[0]) ? 
                       fgallag0x00000_102_q: 
                       fgallag0x00000_103_q;
              fgallag0x00001_52 = 
          (!fgallag_sel[0]) ? 
                       fgallag0x00000_104_q: 
                       fgallag0x00000_105_q;
              fgallag0x00001_53 = 
          (!fgallag_sel[0]) ? 
                       fgallag0x00000_106_q: 
                       fgallag0x00000_107_q;
               fgallag0x00001_54 =  fgallag0x00000_108_q ;
               fgallag0x00001_55 =  fgallag0x00000_110_q ;
              fgallag0x00001_56 = 
          (!fgallag_sel[0]) ? 
                       fgallag0x00000_112_q: 
                       fgallag0x00000_113_q;
               fgallag0x00001_57 =  fgallag0x00000_114_q ;
               fgallag0x00001_58 =  fgallag0x00000_116_q ;
              fgallag0x00001_59 = 
          (!fgallag_sel[0]) ? 
                       fgallag0x00000_118_q: 
                       fgallag0x00000_119_q;
               fgallag0x00001_60 =  fgallag0x00000_120_q ;
               fgallag0x00001_61 =  fgallag0x00000_122_q ;
              fgallag0x00001_62 = 
          (!fgallag_sel[0]) ? 
                       fgallag0x00000_124_q: 
                       fgallag0x00000_125_q;
               fgallag0x00001_63 =  fgallag0x00000_126_q ;
              fgallag0x00001_64 = 
          (!fgallag_sel[0]) ? 
                       fgallag0x00000_128_q: 
                       fgallag0x00000_129_q;
               fgallag0x00001_65 =  fgallag0x00000_130_q ;
               fgallag0x00001_66 =  fgallag0x00000_132_q ;
               fgallag0x00001_67 =  fgallag0x00000_134_q ;
               fgallag0x00001_68 =  fgallag0x00000_136_q ;
               fgallag0x00001_69 =  fgallag0x00000_138_q ;
               fgallag0x00001_70 =  fgallag0x00000_140_q ;
               fgallag0x00001_71 =  fgallag0x00000_142_q ;
              fgallag0x00001_72 = 
          (!fgallag_sel[0]) ? 
                       fgallag0x00000_144_q: 
                       fgallag0x00000_145_q;
               fgallag0x00001_73 =  fgallag0x00000_146_q ;
               fgallag0x00001_74 =  fgallag0x00000_148_q ;
               fgallag0x00001_75 =  fgallag0x00000_150_q ;
               fgallag0x00001_76 =  fgallag0x00000_152_q ;
              fgallag0x00001_77 = 
          (!fgallag_sel[0]) ? 
                       fgallag0x00000_154_q: 
                       fgallag0x00000_155_q;
               fgallag0x00001_78 =  fgallag0x00000_156_q ;
               fgallag0x00001_79 =  fgallag0x00000_158_q ;
              fgallag0x00001_80 = 
          (!fgallag_sel[0]) ? 
                       fgallag0x00000_160_q: 
                       fgallag0x00000_161_q;
               fgallag0x00001_81 =  fgallag0x00000_162_q ;
               fgallag0x00001_82 =  fgallag0x00000_164_q ;
              fgallag0x00001_83 = 
          (!fgallag_sel[0]) ? 
                       fgallag0x00000_166_q: 
                       fgallag0x00000_167_q;
               fgallag0x00001_84 =  fgallag0x00000_168_q ;
               fgallag0x00001_85 =  fgallag0x00000_170_q ;
               fgallag0x00001_86 =  fgallag0x00000_172_q ;
               fgallag0x00001_87 =  fgallag0x00000_174_q ;
               fgallag0x00001_88 =  fgallag0x00000_176_q ;
               fgallag0x00001_89 =  fgallag0x00000_178_q ;
               fgallag0x00001_90 =  fgallag0x00000_180_q ;
               fgallag0x00001_91 =  fgallag0x00000_182_q ;
               fgallag0x00001_92 =  fgallag0x00000_184_q ;
               fgallag0x00001_93 =  fgallag0x00000_186_q ;
               fgallag0x00001_94 =  fgallag0x00000_188_q ;
               fgallag0x00001_95 =  fgallag0x00000_190_q ;
               fgallag0x00001_96 =  fgallag0x00000_192_q ;
               fgallag0x00001_97 =  fgallag0x00000_194_q ;
               fgallag0x00001_98 =  fgallag0x00000_196_q ;
               fgallag0x00001_99 =  fgallag0x00000_198_q ;
               fgallag0x00001_100 =  fgallag0x00000_200_q ;
               fgallag0x00001_101 =  fgallag0x00000_202_q ;
               fgallag0x00001_102 =  fgallag0x00000_204_q ;
               fgallag0x00001_103 =  fgallag0x00000_206_q ;
               fgallag0x00001_104 =  fgallag0x00000_208_q ;
               fgallag0x00001_105 =  fgallag0x00000_210_q ;
               fgallag0x00001_106 =  fgallag0x00000_212_q ;
              fgallag0x00001_107 = 
          (!fgallag_sel[0]) ? 
                       fgallag0x00000_214_q: 
                       fgallag0x00000_215_q;
               fgallag0x00001_108 =  fgallag0x00000_216_q ;
               fgallag0x00001_109 =  fgallag0x00000_218_q ;
               fgallag0x00001_110 =  fgallag0x00000_220_q ;
               fgallag0x00001_111 =  fgallag0x00000_222_q ;
               fgallag0x00001_112 =  fgallag0x00000_224_q ;
               fgallag0x00001_113 =  fgallag0x00000_226_q ;
               fgallag0x00001_114 =  fgallag0x00000_228_q ;
              fgallag0x00001_115 = 
          (!fgallag_sel[0]) ? 
                       fgallag0x00000_230_q: 
                       fgallag0x00000_231_q;
               fgallag0x00001_116 =  fgallag0x00000_232_q ;
               fgallag0x00001_117 =  fgallag0x00000_234_q ;
               fgallag0x00001_118 =  fgallag0x00000_236_q ;
               fgallag0x00001_119 =  fgallag0x00000_238_q ;
               fgallag0x00001_120 =  fgallag0x00000_240_q ;
               fgallag0x00001_121 =  fgallag0x00000_242_q ;
               fgallag0x00001_122 =  fgallag0x00000_244_q ;
               fgallag0x00001_123 =  fgallag0x00000_246_q ;
               fgallag0x00001_124 =  fgallag0x00000_248_q ;
               fgallag0x00001_125 =  fgallag0x00000_250_q ;
              fgallag0x00001_126 = 
          (!fgallag_sel[0]) ? 
                       fgallag0x00000_252_q: 
                       fgallag0x00000_253_q;
               fgallag0x00001_127 =  fgallag0x00000_254_q ;
               fgallag0x00001_128 =  fgallag0x00000_256_q ;
               fgallag0x00001_129 =  fgallag0x00000_258_q ;
               fgallag0x00001_130 =  fgallag0x00000_260_q ;
               fgallag0x00001_131 =  fgallag0x00000_262_q ;
               fgallag0x00001_132 =  fgallag0x00000_264_q ;
               fgallag0x00001_133 =  fgallag0x00000_266_q ;
               fgallag0x00001_134 =  fgallag0x00000_268_q ;
               fgallag0x00001_135 =  fgallag0x00000_270_q ;
               fgallag0x00001_136 =  fgallag0x00000_272_q ;
               fgallag0x00001_137 =  fgallag0x00000_274_q ;
               fgallag0x00001_138 =  fgallag0x00000_276_q ;
               fgallag0x00001_139 =  fgallag0x00000_278_q ;
               fgallag0x00001_140 =  fgallag0x00000_280_q ;
               fgallag0x00001_141 =  fgallag0x00000_282_q ;
              fgallag0x00001_142 = 
          (!fgallag_sel[0]) ? 
                       fgallag0x00000_284_q: 
                       fgallag0x00000_285_q;
               fgallag0x00001_143 =  fgallag0x00000_286_q ;
               fgallag0x00001_144 =  fgallag0x00000_288_q ;
               fgallag0x00001_145 =  fgallag0x00000_290_q ;
               fgallag0x00001_146 =  fgallag0x00000_292_q ;
               fgallag0x00001_147 =  fgallag0x00000_294_q ;
               fgallag0x00001_148 =  fgallag0x00000_296_q ;
               fgallag0x00001_149 =  fgallag0x00000_298_q ;
               fgallag0x00001_150 =  fgallag0x00000_300_q ;
               fgallag0x00001_151 =  fgallag0x00000_302_q ;
               fgallag0x00001_152 =  fgallag0x00000_304_q ;
               fgallag0x00001_153 =  fgallag0x00000_306_q ;
               fgallag0x00001_154 =  fgallag0x00000_308_q ;
               fgallag0x00001_155 =  fgallag0x00000_310_q ;
               fgallag0x00001_156 =  fgallag0x00000_312_q ;
               fgallag0x00001_157 =  fgallag0x00000_314_q ;
               fgallag0x00001_158 =  fgallag0x00000_316_q ;
               fgallag0x00001_159 =  fgallag0x00000_318_q ;
               fgallag0x00001_160 =  fgallag0x00000_320_q ;
               fgallag0x00001_161 =  fgallag0x00000_322_q ;
               fgallag0x00001_162 =  fgallag0x00000_324_q ;
               fgallag0x00001_163 =  fgallag0x00000_326_q ;
               fgallag0x00001_164 =  fgallag0x00000_328_q ;
               fgallag0x00001_165 =  fgallag0x00000_330_q ;
               fgallag0x00001_166 =  fgallag0x00000_332_q ;
               fgallag0x00001_167 =  fgallag0x00000_334_q ;
               fgallag0x00001_168 =  fgallag0x00000_336_q ;
               fgallag0x00001_169 =  fgallag0x00000_338_q ;
               fgallag0x00001_170 =  fgallag0x00000_340_q ;
               fgallag0x00001_171 =  fgallag0x00000_342_q ;
               fgallag0x00001_172 =  fgallag0x00000_344_q ;
               fgallag0x00001_173 =  fgallag0x00000_346_q ;
               fgallag0x00001_174 =  fgallag0x00000_348_q ;
               fgallag0x00001_175 =  fgallag0x00000_350_q ;
               fgallag0x00001_176 =  fgallag0x00000_352_q ;
               fgallag0x00001_177 =  fgallag0x00000_354_q ;
