reg [fgallag_WDTH -1:0] fgallag0x00001_0, fgallag0x00001_0_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_1, fgallag0x00001_1_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_2, fgallag0x00001_2_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_3, fgallag0x00001_3_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_4, fgallag0x00001_4_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_5, fgallag0x00001_5_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_6, fgallag0x00001_6_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_7, fgallag0x00001_7_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_8, fgallag0x00001_8_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_9, fgallag0x00001_9_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_10, fgallag0x00001_10_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_11, fgallag0x00001_11_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_12, fgallag0x00001_12_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_13, fgallag0x00001_13_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_14, fgallag0x00001_14_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_15, fgallag0x00001_15_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_16, fgallag0x00001_16_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_17, fgallag0x00001_17_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_18, fgallag0x00001_18_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_19, fgallag0x00001_19_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_20, fgallag0x00001_20_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_21, fgallag0x00001_21_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_22, fgallag0x00001_22_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_23, fgallag0x00001_23_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_24, fgallag0x00001_24_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_25, fgallag0x00001_25_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_26, fgallag0x00001_26_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_27, fgallag0x00001_27_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_28, fgallag0x00001_28_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_29, fgallag0x00001_29_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_30, fgallag0x00001_30_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_31, fgallag0x00001_31_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_32, fgallag0x00001_32_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_33, fgallag0x00001_33_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_34, fgallag0x00001_34_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_35, fgallag0x00001_35_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_36, fgallag0x00001_36_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_37, fgallag0x00001_37_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_38, fgallag0x00001_38_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_39, fgallag0x00001_39_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_40, fgallag0x00001_40_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_41, fgallag0x00001_41_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_42, fgallag0x00001_42_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_43, fgallag0x00001_43_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_44, fgallag0x00001_44_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_45, fgallag0x00001_45_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_46, fgallag0x00001_46_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_47, fgallag0x00001_47_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_48, fgallag0x00001_48_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_49, fgallag0x00001_49_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_50, fgallag0x00001_50_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_51, fgallag0x00001_51_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_52, fgallag0x00001_52_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_53, fgallag0x00001_53_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_54, fgallag0x00001_54_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_55, fgallag0x00001_55_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_56, fgallag0x00001_56_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_57, fgallag0x00001_57_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_58, fgallag0x00001_58_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_59, fgallag0x00001_59_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_60, fgallag0x00001_60_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_61, fgallag0x00001_61_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_62, fgallag0x00001_62_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_63, fgallag0x00001_63_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_64, fgallag0x00001_64_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_65, fgallag0x00001_65_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_66, fgallag0x00001_66_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_67, fgallag0x00001_67_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_68, fgallag0x00001_68_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_69, fgallag0x00001_69_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_70, fgallag0x00001_70_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_71, fgallag0x00001_71_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_72, fgallag0x00001_72_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_73, fgallag0x00001_73_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_74, fgallag0x00001_74_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_75, fgallag0x00001_75_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_76, fgallag0x00001_76_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_77, fgallag0x00001_77_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_78, fgallag0x00001_78_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_79, fgallag0x00001_79_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_80, fgallag0x00001_80_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_81, fgallag0x00001_81_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_82, fgallag0x00001_82_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_83, fgallag0x00001_83_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_84, fgallag0x00001_84_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_85, fgallag0x00001_85_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_86, fgallag0x00001_86_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_87, fgallag0x00001_87_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_88, fgallag0x00001_88_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_89, fgallag0x00001_89_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_90, fgallag0x00001_90_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_91, fgallag0x00001_91_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_92, fgallag0x00001_92_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_93, fgallag0x00001_93_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_94, fgallag0x00001_94_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_95, fgallag0x00001_95_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_96, fgallag0x00001_96_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_97, fgallag0x00001_97_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_98, fgallag0x00001_98_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_99, fgallag0x00001_99_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_100, fgallag0x00001_100_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_101, fgallag0x00001_101_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_102, fgallag0x00001_102_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_103, fgallag0x00001_103_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_104, fgallag0x00001_104_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_105, fgallag0x00001_105_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_106, fgallag0x00001_106_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_107, fgallag0x00001_107_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_108, fgallag0x00001_108_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_109, fgallag0x00001_109_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_110, fgallag0x00001_110_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_111, fgallag0x00001_111_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_112, fgallag0x00001_112_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_113, fgallag0x00001_113_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_114, fgallag0x00001_114_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_115, fgallag0x00001_115_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_116, fgallag0x00001_116_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_117, fgallag0x00001_117_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_118, fgallag0x00001_118_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_119, fgallag0x00001_119_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_120, fgallag0x00001_120_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_121, fgallag0x00001_121_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_122, fgallag0x00001_122_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_123, fgallag0x00001_123_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_124, fgallag0x00001_124_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_125, fgallag0x00001_125_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_126, fgallag0x00001_126_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_127, fgallag0x00001_127_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_128, fgallag0x00001_128_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_129, fgallag0x00001_129_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_130, fgallag0x00001_130_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_131, fgallag0x00001_131_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_132, fgallag0x00001_132_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_133, fgallag0x00001_133_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_134, fgallag0x00001_134_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_135, fgallag0x00001_135_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_136, fgallag0x00001_136_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_137, fgallag0x00001_137_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_138, fgallag0x00001_138_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_139, fgallag0x00001_139_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_140, fgallag0x00001_140_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_141, fgallag0x00001_141_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_142, fgallag0x00001_142_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_143, fgallag0x00001_143_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_144, fgallag0x00001_144_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_145, fgallag0x00001_145_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_146, fgallag0x00001_146_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_147, fgallag0x00001_147_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_148, fgallag0x00001_148_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_149, fgallag0x00001_149_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_150, fgallag0x00001_150_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_151, fgallag0x00001_151_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_152, fgallag0x00001_152_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_153, fgallag0x00001_153_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_154, fgallag0x00001_154_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_155, fgallag0x00001_155_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_156, fgallag0x00001_156_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_157, fgallag0x00001_157_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_158, fgallag0x00001_158_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_159, fgallag0x00001_159_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_160, fgallag0x00001_160_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_161, fgallag0x00001_161_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_162, fgallag0x00001_162_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_163, fgallag0x00001_163_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_164, fgallag0x00001_164_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_165, fgallag0x00001_165_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_166, fgallag0x00001_166_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_167, fgallag0x00001_167_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_168, fgallag0x00001_168_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_169, fgallag0x00001_169_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_170, fgallag0x00001_170_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_171, fgallag0x00001_171_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_172, fgallag0x00001_172_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_173, fgallag0x00001_173_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_174, fgallag0x00001_174_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_175, fgallag0x00001_175_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_176, fgallag0x00001_176_q;
reg [fgallag_WDTH -1:0] fgallag0x00001_177, fgallag0x00001_177_q;
reg start_d_fgallag0x00001_q ;
always_comb begin
 fgallag0x00001_0_q =  fgallag0x00001_0;
 fgallag0x00001_1_q =  fgallag0x00001_1;
 fgallag0x00001_2_q =  fgallag0x00001_2;
 fgallag0x00001_3_q =  fgallag0x00001_3;
 fgallag0x00001_4_q =  fgallag0x00001_4;
 fgallag0x00001_5_q =  fgallag0x00001_5;
 fgallag0x00001_6_q =  fgallag0x00001_6;
 fgallag0x00001_7_q =  fgallag0x00001_7;
 fgallag0x00001_8_q =  fgallag0x00001_8;
 fgallag0x00001_9_q =  fgallag0x00001_9;
 fgallag0x00001_10_q =  fgallag0x00001_10;
 fgallag0x00001_11_q =  fgallag0x00001_11;
 fgallag0x00001_12_q =  fgallag0x00001_12;
 fgallag0x00001_13_q =  fgallag0x00001_13;
 fgallag0x00001_14_q =  fgallag0x00001_14;
 fgallag0x00001_15_q =  fgallag0x00001_15;
 fgallag0x00001_16_q =  fgallag0x00001_16;
 fgallag0x00001_17_q =  fgallag0x00001_17;
 fgallag0x00001_18_q =  fgallag0x00001_18;
 fgallag0x00001_19_q =  fgallag0x00001_19;
 fgallag0x00001_20_q =  fgallag0x00001_20;
 fgallag0x00001_21_q =  fgallag0x00001_21;
 fgallag0x00001_22_q =  fgallag0x00001_22;
 fgallag0x00001_23_q =  fgallag0x00001_23;
 fgallag0x00001_24_q =  fgallag0x00001_24;
 fgallag0x00001_25_q =  fgallag0x00001_25;
 fgallag0x00001_26_q =  fgallag0x00001_26;
 fgallag0x00001_27_q =  fgallag0x00001_27;
 fgallag0x00001_28_q =  fgallag0x00001_28;
 fgallag0x00001_29_q =  fgallag0x00001_29;
 fgallag0x00001_30_q =  fgallag0x00001_30;
 fgallag0x00001_31_q =  fgallag0x00001_31;
 fgallag0x00001_32_q =  fgallag0x00001_32;
 fgallag0x00001_33_q =  fgallag0x00001_33;
 fgallag0x00001_34_q =  fgallag0x00001_34;
 fgallag0x00001_35_q =  fgallag0x00001_35;
 fgallag0x00001_36_q =  fgallag0x00001_36;
 fgallag0x00001_37_q =  fgallag0x00001_37;
 fgallag0x00001_38_q =  fgallag0x00001_38;
 fgallag0x00001_39_q =  fgallag0x00001_39;
 fgallag0x00001_40_q =  fgallag0x00001_40;
 fgallag0x00001_41_q =  fgallag0x00001_41;
 fgallag0x00001_42_q =  fgallag0x00001_42;
 fgallag0x00001_43_q =  fgallag0x00001_43;
 fgallag0x00001_44_q =  fgallag0x00001_44;
 fgallag0x00001_45_q =  fgallag0x00001_45;
 fgallag0x00001_46_q =  fgallag0x00001_46;
 fgallag0x00001_47_q =  fgallag0x00001_47;
 fgallag0x00001_48_q =  fgallag0x00001_48;
 fgallag0x00001_49_q =  fgallag0x00001_49;
 fgallag0x00001_50_q =  fgallag0x00001_50;
 fgallag0x00001_51_q =  fgallag0x00001_51;
 fgallag0x00001_52_q =  fgallag0x00001_52;
 fgallag0x00001_53_q =  fgallag0x00001_53;
 fgallag0x00001_54_q =  fgallag0x00001_54;
 fgallag0x00001_55_q =  fgallag0x00001_55;
 fgallag0x00001_56_q =  fgallag0x00001_56;
 fgallag0x00001_57_q =  fgallag0x00001_57;
 fgallag0x00001_58_q =  fgallag0x00001_58;
 fgallag0x00001_59_q =  fgallag0x00001_59;
 fgallag0x00001_60_q =  fgallag0x00001_60;
 fgallag0x00001_61_q =  fgallag0x00001_61;
 fgallag0x00001_62_q =  fgallag0x00001_62;
 fgallag0x00001_63_q =  fgallag0x00001_63;
 fgallag0x00001_64_q =  fgallag0x00001_64;
 fgallag0x00001_65_q =  fgallag0x00001_65;
 fgallag0x00001_66_q =  fgallag0x00001_66;
 fgallag0x00001_67_q =  fgallag0x00001_67;
 fgallag0x00001_68_q =  fgallag0x00001_68;
 fgallag0x00001_69_q =  fgallag0x00001_69;
 fgallag0x00001_70_q =  fgallag0x00001_70;
 fgallag0x00001_71_q =  fgallag0x00001_71;
 fgallag0x00001_72_q =  fgallag0x00001_72;
 fgallag0x00001_73_q =  fgallag0x00001_73;
 fgallag0x00001_74_q =  fgallag0x00001_74;
 fgallag0x00001_75_q =  fgallag0x00001_75;
 fgallag0x00001_76_q =  fgallag0x00001_76;
 fgallag0x00001_77_q =  fgallag0x00001_77;
 fgallag0x00001_78_q =  fgallag0x00001_78;
 fgallag0x00001_79_q =  fgallag0x00001_79;
 fgallag0x00001_80_q =  fgallag0x00001_80;
 fgallag0x00001_81_q =  fgallag0x00001_81;
 fgallag0x00001_82_q =  fgallag0x00001_82;
 fgallag0x00001_83_q =  fgallag0x00001_83;
 fgallag0x00001_84_q =  fgallag0x00001_84;
 fgallag0x00001_85_q =  fgallag0x00001_85;
 fgallag0x00001_86_q =  fgallag0x00001_86;
 fgallag0x00001_87_q =  fgallag0x00001_87;
 fgallag0x00001_88_q =  fgallag0x00001_88;
 fgallag0x00001_89_q =  fgallag0x00001_89;
 fgallag0x00001_90_q =  fgallag0x00001_90;
 fgallag0x00001_91_q =  fgallag0x00001_91;
 fgallag0x00001_92_q =  fgallag0x00001_92;
 fgallag0x00001_93_q =  fgallag0x00001_93;
 fgallag0x00001_94_q =  fgallag0x00001_94;
 fgallag0x00001_95_q =  fgallag0x00001_95;
 fgallag0x00001_96_q =  fgallag0x00001_96;
 fgallag0x00001_97_q =  fgallag0x00001_97;
 fgallag0x00001_98_q =  fgallag0x00001_98;
 fgallag0x00001_99_q =  fgallag0x00001_99;
 fgallag0x00001_100_q =  fgallag0x00001_100;
 fgallag0x00001_101_q =  fgallag0x00001_101;
 fgallag0x00001_102_q =  fgallag0x00001_102;
 fgallag0x00001_103_q =  fgallag0x00001_103;
 fgallag0x00001_104_q =  fgallag0x00001_104;
 fgallag0x00001_105_q =  fgallag0x00001_105;
 fgallag0x00001_106_q =  fgallag0x00001_106;
 fgallag0x00001_107_q =  fgallag0x00001_107;
 fgallag0x00001_108_q =  fgallag0x00001_108;
 fgallag0x00001_109_q =  fgallag0x00001_109;
 fgallag0x00001_110_q =  fgallag0x00001_110;
 fgallag0x00001_111_q =  fgallag0x00001_111;
 fgallag0x00001_112_q =  fgallag0x00001_112;
 fgallag0x00001_113_q =  fgallag0x00001_113;
 fgallag0x00001_114_q =  fgallag0x00001_114;
 fgallag0x00001_115_q =  fgallag0x00001_115;
 fgallag0x00001_116_q =  fgallag0x00001_116;
 fgallag0x00001_117_q =  fgallag0x00001_117;
 fgallag0x00001_118_q =  fgallag0x00001_118;
 fgallag0x00001_119_q =  fgallag0x00001_119;
 fgallag0x00001_120_q =  fgallag0x00001_120;
 fgallag0x00001_121_q =  fgallag0x00001_121;
 fgallag0x00001_122_q =  fgallag0x00001_122;
 fgallag0x00001_123_q =  fgallag0x00001_123;
 fgallag0x00001_124_q =  fgallag0x00001_124;
 fgallag0x00001_125_q =  fgallag0x00001_125;
 fgallag0x00001_126_q =  fgallag0x00001_126;
 fgallag0x00001_127_q =  fgallag0x00001_127;
 fgallag0x00001_128_q =  fgallag0x00001_128;
 fgallag0x00001_129_q =  fgallag0x00001_129;
 fgallag0x00001_130_q =  fgallag0x00001_130;
 fgallag0x00001_131_q =  fgallag0x00001_131;
 fgallag0x00001_132_q =  fgallag0x00001_132;
 fgallag0x00001_133_q =  fgallag0x00001_133;
 fgallag0x00001_134_q =  fgallag0x00001_134;
 fgallag0x00001_135_q =  fgallag0x00001_135;
 fgallag0x00001_136_q =  fgallag0x00001_136;
 fgallag0x00001_137_q =  fgallag0x00001_137;
 fgallag0x00001_138_q =  fgallag0x00001_138;
 fgallag0x00001_139_q =  fgallag0x00001_139;
 fgallag0x00001_140_q =  fgallag0x00001_140;
 fgallag0x00001_141_q =  fgallag0x00001_141;
 fgallag0x00001_142_q =  fgallag0x00001_142;
 fgallag0x00001_143_q =  fgallag0x00001_143;
 fgallag0x00001_144_q =  fgallag0x00001_144;
 fgallag0x00001_145_q =  fgallag0x00001_145;
 fgallag0x00001_146_q =  fgallag0x00001_146;
 fgallag0x00001_147_q =  fgallag0x00001_147;
 fgallag0x00001_148_q =  fgallag0x00001_148;
 fgallag0x00001_149_q =  fgallag0x00001_149;
 fgallag0x00001_150_q =  fgallag0x00001_150;
 fgallag0x00001_151_q =  fgallag0x00001_151;
 fgallag0x00001_152_q =  fgallag0x00001_152;
 fgallag0x00001_153_q =  fgallag0x00001_153;
 fgallag0x00001_154_q =  fgallag0x00001_154;
 fgallag0x00001_155_q =  fgallag0x00001_155;
 fgallag0x00001_156_q =  fgallag0x00001_156;
 fgallag0x00001_157_q =  fgallag0x00001_157;
 fgallag0x00001_158_q =  fgallag0x00001_158;
 fgallag0x00001_159_q =  fgallag0x00001_159;
 fgallag0x00001_160_q =  fgallag0x00001_160;
 fgallag0x00001_161_q =  fgallag0x00001_161;
 fgallag0x00001_162_q =  fgallag0x00001_162;
 fgallag0x00001_163_q =  fgallag0x00001_163;
 fgallag0x00001_164_q =  fgallag0x00001_164;
 fgallag0x00001_165_q =  fgallag0x00001_165;
 fgallag0x00001_166_q =  fgallag0x00001_166;
 fgallag0x00001_167_q =  fgallag0x00001_167;
 fgallag0x00001_168_q =  fgallag0x00001_168;
 fgallag0x00001_169_q =  fgallag0x00001_169;
 fgallag0x00001_170_q =  fgallag0x00001_170;
 fgallag0x00001_171_q =  fgallag0x00001_171;
 fgallag0x00001_172_q =  fgallag0x00001_172;
 fgallag0x00001_173_q =  fgallag0x00001_173;
 fgallag0x00001_174_q =  fgallag0x00001_174;
 fgallag0x00001_175_q =  fgallag0x00001_175;
 fgallag0x00001_176_q =  fgallag0x00001_176;
 fgallag0x00001_177_q =  fgallag0x00001_177;
 start_d_fgallag0x00001_q =  start_d_fgallag0x00000_q;
end
