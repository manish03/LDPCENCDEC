              flogtanh0x00007_0 = 
          (!flogtanh_sel[6]) ? 
                       flogtanh0x00006_0_q: 
                       flogtanh0x00006_1_q;
              flogtanh0x00007_1 = 
          (!flogtanh_sel[6]) ? 
                       flogtanh0x00006_2_q: 
                       flogtanh0x00006_3_q;
              flogtanh0x00007_2 = 
          (!flogtanh_sel[6]) ? 
                       flogtanh0x00006_4_q: 
                       flogtanh0x00006_5_q;
               flogtanh0x00007_3 =  0;
