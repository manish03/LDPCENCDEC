parameter fgallag_WDTH = 10 ,
parameter fgallag_MAX = 'h380 ,
parameter fgallag_LIMIT_MAX = 'h800 ,
parameter fgallag_LIMIT = 'h164 ,
parameter fgallag_LEN = 'h164 ,
parameter fgallag_SEL = 9
