`define USE_POWER_PINS
