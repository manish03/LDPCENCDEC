package LDPC_CSR_rtl_pkg;
  localparam int LDPC_ENC_MSG_IN_0_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_0_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_0_BYTE_OFFSET = 13'h0000;
  localparam int LDPC_ENC_MSG_IN_0_MSG_INR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_0_MSG_INR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_0_MSG_INR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_0_MSG_INW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_0_MSG_INW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_0_MSG_INW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_MSG_IN_0_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_MSG_IN_0_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_MSG_IN_0_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_MSG_IN_1_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_1_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_1_BYTE_OFFSET = 13'h0004;
  localparam int LDPC_ENC_MSG_IN_1_MSG_INR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_1_MSG_INR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_1_MSG_INR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_1_MSG_INW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_1_MSG_INW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_1_MSG_INW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_MSG_IN_1_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_MSG_IN_1_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_MSG_IN_1_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_MSG_IN_2_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_2_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_2_BYTE_OFFSET = 13'h0008;
  localparam int LDPC_ENC_MSG_IN_2_MSG_INR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_2_MSG_INR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_2_MSG_INR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_2_MSG_INW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_2_MSG_INW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_2_MSG_INW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_MSG_IN_2_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_MSG_IN_2_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_MSG_IN_2_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_MSG_IN_3_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_3_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_3_BYTE_OFFSET = 13'h000c;
  localparam int LDPC_ENC_MSG_IN_3_MSG_INR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_3_MSG_INR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_3_MSG_INR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_3_MSG_INW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_3_MSG_INW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_3_MSG_INW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_MSG_IN_3_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_MSG_IN_3_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_MSG_IN_3_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_MSG_IN_4_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_4_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_4_BYTE_OFFSET = 13'h0010;
  localparam int LDPC_ENC_MSG_IN_4_MSG_INR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_4_MSG_INR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_4_MSG_INR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_4_MSG_INW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_4_MSG_INW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_4_MSG_INW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_MSG_IN_4_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_MSG_IN_4_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_MSG_IN_4_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_MSG_IN_5_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_5_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_5_BYTE_OFFSET = 13'h0014;
  localparam int LDPC_ENC_MSG_IN_5_MSG_INR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_5_MSG_INR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_5_MSG_INR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_5_MSG_INW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_5_MSG_INW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_5_MSG_INW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_MSG_IN_5_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_MSG_IN_5_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_MSG_IN_5_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_MSG_IN_6_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_6_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_6_BYTE_OFFSET = 13'h0018;
  localparam int LDPC_ENC_MSG_IN_6_MSG_INR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_6_MSG_INR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_6_MSG_INR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_6_MSG_INW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_6_MSG_INW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_6_MSG_INW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_MSG_IN_6_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_MSG_IN_6_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_MSG_IN_6_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_MSG_IN_7_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_7_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_7_BYTE_OFFSET = 13'h001c;
  localparam int LDPC_ENC_MSG_IN_7_MSG_INR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_7_MSG_INR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_7_MSG_INR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_7_MSG_INW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_7_MSG_INW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_7_MSG_INW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_MSG_IN_7_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_MSG_IN_7_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_MSG_IN_7_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_MSG_IN_8_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_8_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_8_BYTE_OFFSET = 13'h0020;
  localparam int LDPC_ENC_MSG_IN_8_MSG_INR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_8_MSG_INR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_8_MSG_INR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_8_MSG_INW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_8_MSG_INW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_8_MSG_INW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_MSG_IN_8_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_MSG_IN_8_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_MSG_IN_8_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_MSG_IN_9_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_9_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_9_BYTE_OFFSET = 13'h0024;
  localparam int LDPC_ENC_MSG_IN_9_MSG_INR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_9_MSG_INR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_9_MSG_INR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_9_MSG_INW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_9_MSG_INW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_9_MSG_INW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_MSG_IN_9_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_MSG_IN_9_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_MSG_IN_9_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_MSG_IN_10_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_10_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_10_BYTE_OFFSET = 13'h0028;
  localparam int LDPC_ENC_MSG_IN_10_MSG_INR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_10_MSG_INR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_10_MSG_INR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_10_MSG_INW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_10_MSG_INW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_10_MSG_INW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_MSG_IN_10_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_MSG_IN_10_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_MSG_IN_10_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_MSG_IN_11_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_11_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_11_BYTE_OFFSET = 13'h002c;
  localparam int LDPC_ENC_MSG_IN_11_MSG_INR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_11_MSG_INR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_11_MSG_INR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_11_MSG_INW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_11_MSG_INW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_11_MSG_INW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_MSG_IN_11_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_MSG_IN_11_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_MSG_IN_11_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_MSG_IN_12_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_12_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_12_BYTE_OFFSET = 13'h0030;
  localparam int LDPC_ENC_MSG_IN_12_MSG_INR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_12_MSG_INR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_12_MSG_INR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_12_MSG_INW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_12_MSG_INW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_12_MSG_INW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_MSG_IN_12_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_MSG_IN_12_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_MSG_IN_12_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_MSG_IN_13_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_13_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_13_BYTE_OFFSET = 13'h0034;
  localparam int LDPC_ENC_MSG_IN_13_MSG_INR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_13_MSG_INR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_13_MSG_INR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_13_MSG_INW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_13_MSG_INW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_13_MSG_INW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_MSG_IN_13_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_MSG_IN_13_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_MSG_IN_13_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_MSG_IN_14_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_14_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_14_BYTE_OFFSET = 13'h0038;
  localparam int LDPC_ENC_MSG_IN_14_MSG_INR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_14_MSG_INR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_14_MSG_INR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_14_MSG_INW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_14_MSG_INW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_14_MSG_INW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_MSG_IN_14_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_MSG_IN_14_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_MSG_IN_14_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_MSG_IN_15_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_15_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_15_BYTE_OFFSET = 13'h003c;
  localparam int LDPC_ENC_MSG_IN_15_MSG_INR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_15_MSG_INR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_15_MSG_INR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_15_MSG_INW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_15_MSG_INW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_15_MSG_INW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_MSG_IN_15_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_MSG_IN_15_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_MSG_IN_15_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_MSG_IN_16_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_16_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_16_BYTE_OFFSET = 13'h0040;
  localparam int LDPC_ENC_MSG_IN_16_MSG_INR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_16_MSG_INR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_16_MSG_INR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_16_MSG_INW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_16_MSG_INW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_16_MSG_INW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_MSG_IN_16_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_MSG_IN_16_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_MSG_IN_16_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_MSG_IN_17_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_17_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_17_BYTE_OFFSET = 13'h0044;
  localparam int LDPC_ENC_MSG_IN_17_MSG_INR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_17_MSG_INR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_17_MSG_INR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_17_MSG_INW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_17_MSG_INW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_17_MSG_INW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_MSG_IN_17_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_MSG_IN_17_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_MSG_IN_17_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_MSG_IN_18_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_18_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_18_BYTE_OFFSET = 13'h0048;
  localparam int LDPC_ENC_MSG_IN_18_MSG_INR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_18_MSG_INR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_18_MSG_INR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_18_MSG_INW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_18_MSG_INW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_18_MSG_INW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_MSG_IN_18_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_MSG_IN_18_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_MSG_IN_18_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_MSG_IN_19_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_19_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_19_BYTE_OFFSET = 13'h004c;
  localparam int LDPC_ENC_MSG_IN_19_MSG_INR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_19_MSG_INR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_19_MSG_INR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_19_MSG_INW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_19_MSG_INW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_19_MSG_INW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_MSG_IN_19_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_MSG_IN_19_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_MSG_IN_19_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_MSG_IN_20_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_20_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_20_BYTE_OFFSET = 13'h0050;
  localparam int LDPC_ENC_MSG_IN_20_MSG_INR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_20_MSG_INR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_20_MSG_INR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_20_MSG_INW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_20_MSG_INW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_20_MSG_INW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_MSG_IN_20_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_MSG_IN_20_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_MSG_IN_20_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_MSG_IN_21_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_21_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_21_BYTE_OFFSET = 13'h0054;
  localparam int LDPC_ENC_MSG_IN_21_MSG_INR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_21_MSG_INR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_21_MSG_INR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_21_MSG_INW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_21_MSG_INW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_21_MSG_INW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_MSG_IN_21_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_MSG_IN_21_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_MSG_IN_21_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_MSG_IN_22_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_22_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_22_BYTE_OFFSET = 13'h0058;
  localparam int LDPC_ENC_MSG_IN_22_MSG_INR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_22_MSG_INR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_22_MSG_INR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_22_MSG_INW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_22_MSG_INW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_22_MSG_INW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_MSG_IN_22_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_MSG_IN_22_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_MSG_IN_22_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_MSG_IN_23_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_23_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_23_BYTE_OFFSET = 13'h005c;
  localparam int LDPC_ENC_MSG_IN_23_MSG_INR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_23_MSG_INR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_23_MSG_INR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_23_MSG_INW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_23_MSG_INW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_23_MSG_INW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_MSG_IN_23_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_MSG_IN_23_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_MSG_IN_23_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_MSG_IN_24_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_24_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_24_BYTE_OFFSET = 13'h0060;
  localparam int LDPC_ENC_MSG_IN_24_MSG_INR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_24_MSG_INR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_24_MSG_INR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_24_MSG_INW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_24_MSG_INW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_24_MSG_INW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_MSG_IN_24_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_MSG_IN_24_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_MSG_IN_24_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_MSG_IN_25_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_25_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_25_BYTE_OFFSET = 13'h0064;
  localparam int LDPC_ENC_MSG_IN_25_MSG_INR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_25_MSG_INR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_25_MSG_INR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_25_MSG_INW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_25_MSG_INW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_25_MSG_INW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_MSG_IN_25_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_MSG_IN_25_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_MSG_IN_25_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_MSG_IN_26_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_26_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_26_BYTE_OFFSET = 13'h0068;
  localparam int LDPC_ENC_MSG_IN_26_MSG_INR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_26_MSG_INR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_26_MSG_INR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_26_MSG_INW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_26_MSG_INW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_26_MSG_INW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_MSG_IN_26_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_MSG_IN_26_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_MSG_IN_26_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_MSG_IN_27_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_27_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_27_BYTE_OFFSET = 13'h006c;
  localparam int LDPC_ENC_MSG_IN_27_MSG_INR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_27_MSG_INR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_27_MSG_INR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_27_MSG_INW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_27_MSG_INW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_27_MSG_INW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_MSG_IN_27_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_MSG_IN_27_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_MSG_IN_27_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_MSG_IN_28_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_28_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_28_BYTE_OFFSET = 13'h0070;
  localparam int LDPC_ENC_MSG_IN_28_MSG_INR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_28_MSG_INR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_28_MSG_INR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_28_MSG_INW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_28_MSG_INW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_28_MSG_INW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_MSG_IN_28_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_MSG_IN_28_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_MSG_IN_28_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_MSG_IN_29_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_29_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_29_BYTE_OFFSET = 13'h0074;
  localparam int LDPC_ENC_MSG_IN_29_MSG_INR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_29_MSG_INR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_29_MSG_INR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_29_MSG_INW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_29_MSG_INW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_29_MSG_INW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_MSG_IN_29_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_MSG_IN_29_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_MSG_IN_29_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_MSG_IN_30_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_30_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_30_BYTE_OFFSET = 13'h0078;
  localparam int LDPC_ENC_MSG_IN_30_MSG_INR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_30_MSG_INR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_30_MSG_INR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_30_MSG_INW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_30_MSG_INW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_30_MSG_INW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_MSG_IN_30_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_MSG_IN_30_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_MSG_IN_30_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_MSG_IN_31_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_31_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_31_BYTE_OFFSET = 13'h007c;
  localparam int LDPC_ENC_MSG_IN_31_MSG_INR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_31_MSG_INR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_31_MSG_INR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_31_MSG_INW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_31_MSG_INW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_31_MSG_INW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_MSG_IN_31_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_MSG_IN_31_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_MSG_IN_31_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_MSG_IN_32_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_32_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_32_BYTE_OFFSET = 13'h0080;
  localparam int LDPC_ENC_MSG_IN_32_MSG_INR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_32_MSG_INR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_32_MSG_INR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_32_MSG_INW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_32_MSG_INW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_32_MSG_INW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_MSG_IN_32_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_MSG_IN_32_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_MSG_IN_32_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_MSG_IN_33_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_33_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_33_BYTE_OFFSET = 13'h0084;
  localparam int LDPC_ENC_MSG_IN_33_MSG_INR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_33_MSG_INR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_33_MSG_INR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_33_MSG_INW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_33_MSG_INW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_33_MSG_INW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_MSG_IN_33_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_MSG_IN_33_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_MSG_IN_33_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_MSG_IN_34_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_34_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_34_BYTE_OFFSET = 13'h0088;
  localparam int LDPC_ENC_MSG_IN_34_MSG_INR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_34_MSG_INR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_34_MSG_INR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_34_MSG_INW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_34_MSG_INW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_34_MSG_INW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_MSG_IN_34_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_MSG_IN_34_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_MSG_IN_34_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_MSG_IN_35_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_35_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_35_BYTE_OFFSET = 13'h008c;
  localparam int LDPC_ENC_MSG_IN_35_MSG_INR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_35_MSG_INR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_35_MSG_INR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_35_MSG_INW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_35_MSG_INW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_35_MSG_INW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_MSG_IN_35_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_MSG_IN_35_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_MSG_IN_35_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_MSG_IN_36_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_36_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_36_BYTE_OFFSET = 13'h0090;
  localparam int LDPC_ENC_MSG_IN_36_MSG_INR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_36_MSG_INR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_36_MSG_INR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_36_MSG_INW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_36_MSG_INW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_36_MSG_INW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_MSG_IN_36_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_MSG_IN_36_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_MSG_IN_36_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_MSG_IN_37_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_37_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_37_BYTE_OFFSET = 13'h0094;
  localparam int LDPC_ENC_MSG_IN_37_MSG_INR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_37_MSG_INR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_37_MSG_INR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_37_MSG_INW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_37_MSG_INW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_37_MSG_INW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_MSG_IN_37_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_MSG_IN_37_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_MSG_IN_37_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_MSG_IN_38_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_38_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_38_BYTE_OFFSET = 13'h0098;
  localparam int LDPC_ENC_MSG_IN_38_MSG_INR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_38_MSG_INR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_38_MSG_INR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_38_MSG_INW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_38_MSG_INW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_38_MSG_INW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_MSG_IN_38_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_MSG_IN_38_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_MSG_IN_38_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_MSG_IN_39_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_39_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_39_BYTE_OFFSET = 13'h009c;
  localparam int LDPC_ENC_MSG_IN_39_MSG_INR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_39_MSG_INR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_39_MSG_INR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_39_MSG_INW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_39_MSG_INW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_39_MSG_INW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_MSG_IN_39_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_MSG_IN_39_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_MSG_IN_39_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_0_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_0_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_0_BYTE_OFFSET = 13'h00a0;
  localparam int LDPC_ENC_CODEWRD_0_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_0_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_0_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_0_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_0_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_0_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_0_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_0_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_0_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_1_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_1_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_1_BYTE_OFFSET = 13'h00a4;
  localparam int LDPC_ENC_CODEWRD_1_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_1_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_1_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_1_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_1_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_1_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_1_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_1_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_1_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_2_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_2_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_2_BYTE_OFFSET = 13'h00a8;
  localparam int LDPC_ENC_CODEWRD_2_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_2_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_2_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_2_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_2_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_2_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_2_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_2_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_2_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_3_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_3_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_3_BYTE_OFFSET = 13'h00ac;
  localparam int LDPC_ENC_CODEWRD_3_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_3_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_3_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_3_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_3_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_3_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_3_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_3_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_3_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_4_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_4_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_4_BYTE_OFFSET = 13'h00b0;
  localparam int LDPC_ENC_CODEWRD_4_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_4_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_4_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_4_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_4_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_4_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_4_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_4_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_4_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_5_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_5_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_5_BYTE_OFFSET = 13'h00b4;
  localparam int LDPC_ENC_CODEWRD_5_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_5_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_5_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_5_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_5_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_5_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_5_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_5_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_5_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_6_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_6_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_6_BYTE_OFFSET = 13'h00b8;
  localparam int LDPC_ENC_CODEWRD_6_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_6_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_6_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_6_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_6_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_6_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_6_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_6_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_6_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_7_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_7_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_7_BYTE_OFFSET = 13'h00bc;
  localparam int LDPC_ENC_CODEWRD_7_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_7_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_7_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_7_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_7_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_7_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_7_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_7_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_7_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_8_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_8_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_8_BYTE_OFFSET = 13'h00c0;
  localparam int LDPC_ENC_CODEWRD_8_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_8_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_8_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_8_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_8_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_8_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_8_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_8_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_8_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_9_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_9_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_9_BYTE_OFFSET = 13'h00c4;
  localparam int LDPC_ENC_CODEWRD_9_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_9_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_9_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_9_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_9_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_9_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_9_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_9_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_9_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_10_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_10_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_10_BYTE_OFFSET = 13'h00c8;
  localparam int LDPC_ENC_CODEWRD_10_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_10_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_10_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_10_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_10_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_10_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_10_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_10_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_10_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_11_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_11_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_11_BYTE_OFFSET = 13'h00cc;
  localparam int LDPC_ENC_CODEWRD_11_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_11_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_11_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_11_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_11_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_11_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_11_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_11_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_11_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_12_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_12_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_12_BYTE_OFFSET = 13'h00d0;
  localparam int LDPC_ENC_CODEWRD_12_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_12_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_12_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_12_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_12_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_12_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_12_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_12_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_12_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_13_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_13_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_13_BYTE_OFFSET = 13'h00d4;
  localparam int LDPC_ENC_CODEWRD_13_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_13_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_13_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_13_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_13_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_13_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_13_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_13_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_13_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_14_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_14_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_14_BYTE_OFFSET = 13'h00d8;
  localparam int LDPC_ENC_CODEWRD_14_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_14_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_14_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_14_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_14_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_14_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_14_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_14_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_14_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_15_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_15_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_15_BYTE_OFFSET = 13'h00dc;
  localparam int LDPC_ENC_CODEWRD_15_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_15_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_15_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_15_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_15_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_15_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_15_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_15_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_15_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_16_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_16_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_16_BYTE_OFFSET = 13'h00e0;
  localparam int LDPC_ENC_CODEWRD_16_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_16_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_16_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_16_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_16_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_16_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_16_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_16_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_16_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_17_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_17_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_17_BYTE_OFFSET = 13'h00e4;
  localparam int LDPC_ENC_CODEWRD_17_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_17_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_17_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_17_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_17_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_17_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_17_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_17_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_17_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_18_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_18_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_18_BYTE_OFFSET = 13'h00e8;
  localparam int LDPC_ENC_CODEWRD_18_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_18_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_18_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_18_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_18_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_18_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_18_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_18_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_18_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_19_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_19_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_19_BYTE_OFFSET = 13'h00ec;
  localparam int LDPC_ENC_CODEWRD_19_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_19_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_19_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_19_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_19_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_19_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_19_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_19_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_19_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_20_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_20_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_20_BYTE_OFFSET = 13'h00f0;
  localparam int LDPC_ENC_CODEWRD_20_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_20_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_20_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_20_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_20_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_20_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_20_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_20_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_20_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_21_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_21_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_21_BYTE_OFFSET = 13'h00f4;
  localparam int LDPC_ENC_CODEWRD_21_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_21_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_21_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_21_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_21_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_21_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_21_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_21_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_21_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_22_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_22_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_22_BYTE_OFFSET = 13'h00f8;
  localparam int LDPC_ENC_CODEWRD_22_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_22_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_22_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_22_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_22_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_22_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_22_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_22_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_22_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_23_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_23_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_23_BYTE_OFFSET = 13'h00fc;
  localparam int LDPC_ENC_CODEWRD_23_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_23_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_23_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_23_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_23_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_23_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_23_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_23_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_23_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_24_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_24_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_24_BYTE_OFFSET = 13'h0100;
  localparam int LDPC_ENC_CODEWRD_24_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_24_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_24_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_24_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_24_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_24_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_24_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_24_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_24_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_25_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_25_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_25_BYTE_OFFSET = 13'h0104;
  localparam int LDPC_ENC_CODEWRD_25_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_25_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_25_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_25_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_25_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_25_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_25_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_25_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_25_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_26_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_26_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_26_BYTE_OFFSET = 13'h0108;
  localparam int LDPC_ENC_CODEWRD_26_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_26_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_26_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_26_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_26_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_26_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_26_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_26_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_26_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_27_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_27_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_27_BYTE_OFFSET = 13'h010c;
  localparam int LDPC_ENC_CODEWRD_27_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_27_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_27_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_27_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_27_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_27_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_27_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_27_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_27_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_28_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_28_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_28_BYTE_OFFSET = 13'h0110;
  localparam int LDPC_ENC_CODEWRD_28_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_28_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_28_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_28_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_28_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_28_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_28_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_28_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_28_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_29_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_29_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_29_BYTE_OFFSET = 13'h0114;
  localparam int LDPC_ENC_CODEWRD_29_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_29_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_29_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_29_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_29_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_29_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_29_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_29_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_29_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_30_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_30_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_30_BYTE_OFFSET = 13'h0118;
  localparam int LDPC_ENC_CODEWRD_30_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_30_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_30_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_30_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_30_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_30_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_30_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_30_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_30_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_31_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_31_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_31_BYTE_OFFSET = 13'h011c;
  localparam int LDPC_ENC_CODEWRD_31_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_31_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_31_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_31_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_31_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_31_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_31_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_31_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_31_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_32_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_32_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_32_BYTE_OFFSET = 13'h0120;
  localparam int LDPC_ENC_CODEWRD_32_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_32_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_32_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_32_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_32_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_32_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_32_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_32_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_32_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_33_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_33_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_33_BYTE_OFFSET = 13'h0124;
  localparam int LDPC_ENC_CODEWRD_33_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_33_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_33_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_33_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_33_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_33_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_33_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_33_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_33_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_34_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_34_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_34_BYTE_OFFSET = 13'h0128;
  localparam int LDPC_ENC_CODEWRD_34_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_34_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_34_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_34_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_34_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_34_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_34_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_34_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_34_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_35_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_35_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_35_BYTE_OFFSET = 13'h012c;
  localparam int LDPC_ENC_CODEWRD_35_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_35_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_35_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_35_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_35_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_35_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_35_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_35_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_35_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_36_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_36_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_36_BYTE_OFFSET = 13'h0130;
  localparam int LDPC_ENC_CODEWRD_36_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_36_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_36_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_36_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_36_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_36_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_36_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_36_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_36_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_37_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_37_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_37_BYTE_OFFSET = 13'h0134;
  localparam int LDPC_ENC_CODEWRD_37_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_37_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_37_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_37_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_37_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_37_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_37_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_37_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_37_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_38_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_38_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_38_BYTE_OFFSET = 13'h0138;
  localparam int LDPC_ENC_CODEWRD_38_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_38_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_38_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_38_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_38_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_38_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_38_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_38_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_38_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_39_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_39_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_39_BYTE_OFFSET = 13'h013c;
  localparam int LDPC_ENC_CODEWRD_39_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_39_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_39_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_39_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_39_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_39_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_39_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_39_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_39_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_40_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_40_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_40_BYTE_OFFSET = 13'h0140;
  localparam int LDPC_ENC_CODEWRD_40_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_40_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_40_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_40_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_40_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_40_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_40_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_40_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_40_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_41_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_41_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_41_BYTE_OFFSET = 13'h0144;
  localparam int LDPC_ENC_CODEWRD_41_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_41_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_41_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_41_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_41_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_41_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_41_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_41_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_41_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_42_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_42_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_42_BYTE_OFFSET = 13'h0148;
  localparam int LDPC_ENC_CODEWRD_42_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_42_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_42_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_42_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_42_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_42_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_42_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_42_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_42_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_43_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_43_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_43_BYTE_OFFSET = 13'h014c;
  localparam int LDPC_ENC_CODEWRD_43_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_43_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_43_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_43_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_43_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_43_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_43_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_43_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_43_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_44_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_44_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_44_BYTE_OFFSET = 13'h0150;
  localparam int LDPC_ENC_CODEWRD_44_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_44_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_44_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_44_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_44_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_44_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_44_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_44_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_44_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_45_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_45_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_45_BYTE_OFFSET = 13'h0154;
  localparam int LDPC_ENC_CODEWRD_45_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_45_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_45_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_45_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_45_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_45_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_45_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_45_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_45_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_46_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_46_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_46_BYTE_OFFSET = 13'h0158;
  localparam int LDPC_ENC_CODEWRD_46_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_46_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_46_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_46_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_46_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_46_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_46_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_46_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_46_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_47_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_47_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_47_BYTE_OFFSET = 13'h015c;
  localparam int LDPC_ENC_CODEWRD_47_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_47_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_47_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_47_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_47_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_47_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_47_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_47_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_47_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_48_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_48_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_48_BYTE_OFFSET = 13'h0160;
  localparam int LDPC_ENC_CODEWRD_48_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_48_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_48_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_48_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_48_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_48_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_48_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_48_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_48_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_49_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_49_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_49_BYTE_OFFSET = 13'h0164;
  localparam int LDPC_ENC_CODEWRD_49_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_49_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_49_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_49_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_49_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_49_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_49_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_49_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_49_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_50_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_50_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_50_BYTE_OFFSET = 13'h0168;
  localparam int LDPC_ENC_CODEWRD_50_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_50_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_50_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_50_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_50_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_50_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_50_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_50_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_50_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_51_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_51_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_51_BYTE_OFFSET = 13'h016c;
  localparam int LDPC_ENC_CODEWRD_51_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_51_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_51_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_51_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_51_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_51_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_51_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_51_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_51_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_52_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_52_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_52_BYTE_OFFSET = 13'h0170;
  localparam int LDPC_ENC_CODEWRD_52_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_52_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_52_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_52_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_52_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_52_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_52_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_52_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_52_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_53_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_53_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_53_BYTE_OFFSET = 13'h0174;
  localparam int LDPC_ENC_CODEWRD_53_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_53_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_53_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_53_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_53_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_53_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_53_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_53_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_53_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_54_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_54_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_54_BYTE_OFFSET = 13'h0178;
  localparam int LDPC_ENC_CODEWRD_54_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_54_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_54_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_54_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_54_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_54_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_54_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_54_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_54_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_55_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_55_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_55_BYTE_OFFSET = 13'h017c;
  localparam int LDPC_ENC_CODEWRD_55_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_55_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_55_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_55_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_55_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_55_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_55_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_55_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_55_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_56_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_56_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_56_BYTE_OFFSET = 13'h0180;
  localparam int LDPC_ENC_CODEWRD_56_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_56_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_56_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_56_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_56_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_56_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_56_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_56_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_56_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_57_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_57_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_57_BYTE_OFFSET = 13'h0184;
  localparam int LDPC_ENC_CODEWRD_57_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_57_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_57_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_57_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_57_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_57_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_57_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_57_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_57_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_58_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_58_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_58_BYTE_OFFSET = 13'h0188;
  localparam int LDPC_ENC_CODEWRD_58_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_58_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_58_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_58_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_58_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_58_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_58_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_58_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_58_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_59_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_59_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_59_BYTE_OFFSET = 13'h018c;
  localparam int LDPC_ENC_CODEWRD_59_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_59_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_59_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_59_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_59_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_59_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_59_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_59_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_59_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_60_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_60_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_60_BYTE_OFFSET = 13'h0190;
  localparam int LDPC_ENC_CODEWRD_60_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_60_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_60_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_60_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_60_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_60_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_60_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_60_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_60_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_61_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_61_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_61_BYTE_OFFSET = 13'h0194;
  localparam int LDPC_ENC_CODEWRD_61_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_61_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_61_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_61_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_61_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_61_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_61_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_61_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_61_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_62_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_62_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_62_BYTE_OFFSET = 13'h0198;
  localparam int LDPC_ENC_CODEWRD_62_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_62_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_62_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_62_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_62_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_62_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_62_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_62_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_62_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_63_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_63_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_63_BYTE_OFFSET = 13'h019c;
  localparam int LDPC_ENC_CODEWRD_63_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_63_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_63_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_63_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_63_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_63_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_63_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_63_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_63_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_64_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_64_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_64_BYTE_OFFSET = 13'h01a0;
  localparam int LDPC_ENC_CODEWRD_64_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_64_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_64_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_64_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_64_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_64_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_64_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_64_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_64_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_65_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_65_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_65_BYTE_OFFSET = 13'h01a4;
  localparam int LDPC_ENC_CODEWRD_65_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_65_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_65_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_65_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_65_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_65_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_65_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_65_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_65_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_66_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_66_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_66_BYTE_OFFSET = 13'h01a8;
  localparam int LDPC_ENC_CODEWRD_66_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_66_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_66_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_66_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_66_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_66_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_66_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_66_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_66_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_67_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_67_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_67_BYTE_OFFSET = 13'h01ac;
  localparam int LDPC_ENC_CODEWRD_67_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_67_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_67_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_67_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_67_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_67_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_67_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_67_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_67_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_68_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_68_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_68_BYTE_OFFSET = 13'h01b0;
  localparam int LDPC_ENC_CODEWRD_68_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_68_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_68_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_68_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_68_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_68_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_68_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_68_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_68_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_69_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_69_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_69_BYTE_OFFSET = 13'h01b4;
  localparam int LDPC_ENC_CODEWRD_69_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_69_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_69_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_69_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_69_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_69_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_69_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_69_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_69_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_70_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_70_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_70_BYTE_OFFSET = 13'h01b8;
  localparam int LDPC_ENC_CODEWRD_70_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_70_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_70_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_70_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_70_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_70_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_70_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_70_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_70_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_71_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_71_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_71_BYTE_OFFSET = 13'h01bc;
  localparam int LDPC_ENC_CODEWRD_71_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_71_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_71_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_71_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_71_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_71_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_71_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_71_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_71_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_72_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_72_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_72_BYTE_OFFSET = 13'h01c0;
  localparam int LDPC_ENC_CODEWRD_72_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_72_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_72_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_72_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_72_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_72_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_72_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_72_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_72_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_73_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_73_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_73_BYTE_OFFSET = 13'h01c4;
  localparam int LDPC_ENC_CODEWRD_73_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_73_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_73_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_73_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_73_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_73_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_73_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_73_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_73_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_74_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_74_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_74_BYTE_OFFSET = 13'h01c8;
  localparam int LDPC_ENC_CODEWRD_74_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_74_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_74_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_74_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_74_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_74_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_74_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_74_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_74_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_75_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_75_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_75_BYTE_OFFSET = 13'h01cc;
  localparam int LDPC_ENC_CODEWRD_75_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_75_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_75_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_75_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_75_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_75_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_75_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_75_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_75_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_76_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_76_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_76_BYTE_OFFSET = 13'h01d0;
  localparam int LDPC_ENC_CODEWRD_76_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_76_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_76_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_76_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_76_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_76_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_76_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_76_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_76_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_77_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_77_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_77_BYTE_OFFSET = 13'h01d4;
  localparam int LDPC_ENC_CODEWRD_77_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_77_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_77_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_77_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_77_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_77_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_77_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_77_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_77_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_78_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_78_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_78_BYTE_OFFSET = 13'h01d8;
  localparam int LDPC_ENC_CODEWRD_78_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_78_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_78_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_78_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_78_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_78_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_78_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_78_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_78_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_79_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_79_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_79_BYTE_OFFSET = 13'h01dc;
  localparam int LDPC_ENC_CODEWRD_79_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_79_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_79_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_79_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_79_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_79_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_79_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_79_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_79_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_80_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_80_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_80_BYTE_OFFSET = 13'h01e0;
  localparam int LDPC_ENC_CODEWRD_80_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_80_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_80_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_80_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_80_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_80_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_80_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_80_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_80_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_81_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_81_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_81_BYTE_OFFSET = 13'h01e4;
  localparam int LDPC_ENC_CODEWRD_81_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_81_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_81_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_81_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_81_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_81_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_81_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_81_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_81_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_82_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_82_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_82_BYTE_OFFSET = 13'h01e8;
  localparam int LDPC_ENC_CODEWRD_82_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_82_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_82_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_82_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_82_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_82_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_82_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_82_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_82_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_83_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_83_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_83_BYTE_OFFSET = 13'h01ec;
  localparam int LDPC_ENC_CODEWRD_83_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_83_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_83_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_83_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_83_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_83_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_83_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_83_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_83_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_84_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_84_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_84_BYTE_OFFSET = 13'h01f0;
  localparam int LDPC_ENC_CODEWRD_84_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_84_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_84_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_84_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_84_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_84_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_84_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_84_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_84_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_85_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_85_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_85_BYTE_OFFSET = 13'h01f4;
  localparam int LDPC_ENC_CODEWRD_85_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_85_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_85_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_85_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_85_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_85_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_85_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_85_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_85_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_86_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_86_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_86_BYTE_OFFSET = 13'h01f8;
  localparam int LDPC_ENC_CODEWRD_86_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_86_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_86_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_86_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_86_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_86_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_86_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_86_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_86_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_87_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_87_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_87_BYTE_OFFSET = 13'h01fc;
  localparam int LDPC_ENC_CODEWRD_87_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_87_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_87_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_87_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_87_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_87_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_87_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_87_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_87_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_88_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_88_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_88_BYTE_OFFSET = 13'h0200;
  localparam int LDPC_ENC_CODEWRD_88_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_88_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_88_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_88_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_88_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_88_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_88_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_88_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_88_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_89_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_89_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_89_BYTE_OFFSET = 13'h0204;
  localparam int LDPC_ENC_CODEWRD_89_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_89_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_89_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_89_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_89_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_89_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_89_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_89_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_89_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_90_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_90_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_90_BYTE_OFFSET = 13'h0208;
  localparam int LDPC_ENC_CODEWRD_90_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_90_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_90_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_90_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_90_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_90_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_90_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_90_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_90_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_91_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_91_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_91_BYTE_OFFSET = 13'h020c;
  localparam int LDPC_ENC_CODEWRD_91_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_91_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_91_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_91_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_91_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_91_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_91_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_91_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_91_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_92_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_92_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_92_BYTE_OFFSET = 13'h0210;
  localparam int LDPC_ENC_CODEWRD_92_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_92_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_92_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_92_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_92_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_92_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_92_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_92_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_92_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_93_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_93_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_93_BYTE_OFFSET = 13'h0214;
  localparam int LDPC_ENC_CODEWRD_93_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_93_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_93_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_93_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_93_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_93_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_93_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_93_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_93_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_94_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_94_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_94_BYTE_OFFSET = 13'h0218;
  localparam int LDPC_ENC_CODEWRD_94_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_94_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_94_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_94_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_94_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_94_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_94_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_94_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_94_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_95_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_95_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_95_BYTE_OFFSET = 13'h021c;
  localparam int LDPC_ENC_CODEWRD_95_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_95_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_95_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_95_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_95_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_95_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_95_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_95_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_95_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_96_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_96_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_96_BYTE_OFFSET = 13'h0220;
  localparam int LDPC_ENC_CODEWRD_96_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_96_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_96_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_96_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_96_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_96_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_96_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_96_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_96_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_97_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_97_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_97_BYTE_OFFSET = 13'h0224;
  localparam int LDPC_ENC_CODEWRD_97_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_97_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_97_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_97_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_97_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_97_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_97_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_97_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_97_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_98_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_98_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_98_BYTE_OFFSET = 13'h0228;
  localparam int LDPC_ENC_CODEWRD_98_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_98_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_98_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_98_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_98_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_98_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_98_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_98_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_98_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_99_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_99_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_99_BYTE_OFFSET = 13'h022c;
  localparam int LDPC_ENC_CODEWRD_99_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_99_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_99_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_99_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_99_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_99_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_99_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_99_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_99_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_100_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_100_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_100_BYTE_OFFSET = 13'h0230;
  localparam int LDPC_ENC_CODEWRD_100_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_100_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_100_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_100_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_100_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_100_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_100_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_100_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_100_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_101_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_101_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_101_BYTE_OFFSET = 13'h0234;
  localparam int LDPC_ENC_CODEWRD_101_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_101_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_101_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_101_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_101_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_101_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_101_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_101_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_101_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_102_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_102_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_102_BYTE_OFFSET = 13'h0238;
  localparam int LDPC_ENC_CODEWRD_102_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_102_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_102_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_102_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_102_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_102_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_102_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_102_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_102_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_103_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_103_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_103_BYTE_OFFSET = 13'h023c;
  localparam int LDPC_ENC_CODEWRD_103_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_103_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_103_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_103_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_103_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_103_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_103_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_103_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_103_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_104_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_104_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_104_BYTE_OFFSET = 13'h0240;
  localparam int LDPC_ENC_CODEWRD_104_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_104_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_104_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_104_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_104_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_104_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_104_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_104_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_104_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_105_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_105_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_105_BYTE_OFFSET = 13'h0244;
  localparam int LDPC_ENC_CODEWRD_105_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_105_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_105_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_105_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_105_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_105_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_105_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_105_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_105_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_106_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_106_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_106_BYTE_OFFSET = 13'h0248;
  localparam int LDPC_ENC_CODEWRD_106_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_106_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_106_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_106_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_106_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_106_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_106_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_106_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_106_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_107_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_107_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_107_BYTE_OFFSET = 13'h024c;
  localparam int LDPC_ENC_CODEWRD_107_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_107_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_107_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_107_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_107_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_107_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_107_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_107_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_107_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_108_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_108_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_108_BYTE_OFFSET = 13'h0250;
  localparam int LDPC_ENC_CODEWRD_108_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_108_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_108_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_108_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_108_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_108_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_108_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_108_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_108_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_109_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_109_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_109_BYTE_OFFSET = 13'h0254;
  localparam int LDPC_ENC_CODEWRD_109_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_109_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_109_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_109_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_109_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_109_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_109_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_109_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_109_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_110_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_110_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_110_BYTE_OFFSET = 13'h0258;
  localparam int LDPC_ENC_CODEWRD_110_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_110_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_110_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_110_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_110_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_110_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_110_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_110_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_110_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_111_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_111_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_111_BYTE_OFFSET = 13'h025c;
  localparam int LDPC_ENC_CODEWRD_111_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_111_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_111_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_111_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_111_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_111_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_111_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_111_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_111_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_112_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_112_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_112_BYTE_OFFSET = 13'h0260;
  localparam int LDPC_ENC_CODEWRD_112_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_112_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_112_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_112_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_112_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_112_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_112_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_112_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_112_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_113_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_113_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_113_BYTE_OFFSET = 13'h0264;
  localparam int LDPC_ENC_CODEWRD_113_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_113_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_113_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_113_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_113_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_113_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_113_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_113_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_113_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_114_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_114_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_114_BYTE_OFFSET = 13'h0268;
  localparam int LDPC_ENC_CODEWRD_114_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_114_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_114_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_114_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_114_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_114_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_114_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_114_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_114_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_115_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_115_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_115_BYTE_OFFSET = 13'h026c;
  localparam int LDPC_ENC_CODEWRD_115_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_115_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_115_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_115_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_115_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_115_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_115_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_115_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_115_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_116_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_116_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_116_BYTE_OFFSET = 13'h0270;
  localparam int LDPC_ENC_CODEWRD_116_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_116_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_116_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_116_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_116_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_116_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_116_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_116_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_116_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_117_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_117_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_117_BYTE_OFFSET = 13'h0274;
  localparam int LDPC_ENC_CODEWRD_117_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_117_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_117_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_117_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_117_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_117_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_117_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_117_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_117_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_118_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_118_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_118_BYTE_OFFSET = 13'h0278;
  localparam int LDPC_ENC_CODEWRD_118_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_118_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_118_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_118_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_118_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_118_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_118_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_118_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_118_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_119_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_119_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_119_BYTE_OFFSET = 13'h027c;
  localparam int LDPC_ENC_CODEWRD_119_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_119_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_119_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_119_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_119_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_119_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_119_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_119_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_119_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_120_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_120_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_120_BYTE_OFFSET = 13'h0280;
  localparam int LDPC_ENC_CODEWRD_120_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_120_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_120_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_120_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_120_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_120_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_120_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_120_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_120_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_121_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_121_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_121_BYTE_OFFSET = 13'h0284;
  localparam int LDPC_ENC_CODEWRD_121_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_121_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_121_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_121_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_121_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_121_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_121_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_121_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_121_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_122_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_122_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_122_BYTE_OFFSET = 13'h0288;
  localparam int LDPC_ENC_CODEWRD_122_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_122_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_122_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_122_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_122_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_122_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_122_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_122_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_122_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_123_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_123_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_123_BYTE_OFFSET = 13'h028c;
  localparam int LDPC_ENC_CODEWRD_123_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_123_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_123_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_123_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_123_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_123_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_123_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_123_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_123_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_124_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_124_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_124_BYTE_OFFSET = 13'h0290;
  localparam int LDPC_ENC_CODEWRD_124_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_124_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_124_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_124_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_124_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_124_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_124_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_124_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_124_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_125_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_125_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_125_BYTE_OFFSET = 13'h0294;
  localparam int LDPC_ENC_CODEWRD_125_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_125_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_125_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_125_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_125_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_125_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_125_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_125_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_125_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_126_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_126_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_126_BYTE_OFFSET = 13'h0298;
  localparam int LDPC_ENC_CODEWRD_126_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_126_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_126_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_126_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_126_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_126_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_126_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_126_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_126_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_127_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_127_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_127_BYTE_OFFSET = 13'h029c;
  localparam int LDPC_ENC_CODEWRD_127_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_127_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_127_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_127_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_127_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_127_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_127_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_127_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_127_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_128_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_128_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_128_BYTE_OFFSET = 13'h02a0;
  localparam int LDPC_ENC_CODEWRD_128_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_128_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_128_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_128_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_128_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_128_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_128_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_128_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_128_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_129_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_129_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_129_BYTE_OFFSET = 13'h02a4;
  localparam int LDPC_ENC_CODEWRD_129_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_129_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_129_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_129_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_129_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_129_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_129_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_129_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_129_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_130_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_130_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_130_BYTE_OFFSET = 13'h02a8;
  localparam int LDPC_ENC_CODEWRD_130_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_130_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_130_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_130_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_130_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_130_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_130_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_130_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_130_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_131_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_131_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_131_BYTE_OFFSET = 13'h02ac;
  localparam int LDPC_ENC_CODEWRD_131_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_131_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_131_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_131_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_131_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_131_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_131_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_131_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_131_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_132_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_132_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_132_BYTE_OFFSET = 13'h02b0;
  localparam int LDPC_ENC_CODEWRD_132_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_132_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_132_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_132_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_132_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_132_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_132_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_132_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_132_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_133_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_133_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_133_BYTE_OFFSET = 13'h02b4;
  localparam int LDPC_ENC_CODEWRD_133_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_133_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_133_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_133_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_133_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_133_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_133_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_133_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_133_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_134_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_134_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_134_BYTE_OFFSET = 13'h02b8;
  localparam int LDPC_ENC_CODEWRD_134_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_134_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_134_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_134_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_134_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_134_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_134_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_134_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_134_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_135_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_135_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_135_BYTE_OFFSET = 13'h02bc;
  localparam int LDPC_ENC_CODEWRD_135_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_135_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_135_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_135_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_135_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_135_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_135_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_135_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_135_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_136_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_136_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_136_BYTE_OFFSET = 13'h02c0;
  localparam int LDPC_ENC_CODEWRD_136_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_136_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_136_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_136_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_136_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_136_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_136_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_136_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_136_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_137_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_137_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_137_BYTE_OFFSET = 13'h02c4;
  localparam int LDPC_ENC_CODEWRD_137_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_137_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_137_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_137_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_137_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_137_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_137_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_137_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_137_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_138_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_138_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_138_BYTE_OFFSET = 13'h02c8;
  localparam int LDPC_ENC_CODEWRD_138_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_138_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_138_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_138_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_138_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_138_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_138_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_138_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_138_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_139_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_139_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_139_BYTE_OFFSET = 13'h02cc;
  localparam int LDPC_ENC_CODEWRD_139_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_139_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_139_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_139_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_139_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_139_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_139_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_139_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_139_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_140_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_140_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_140_BYTE_OFFSET = 13'h02d0;
  localparam int LDPC_ENC_CODEWRD_140_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_140_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_140_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_140_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_140_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_140_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_140_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_140_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_140_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_141_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_141_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_141_BYTE_OFFSET = 13'h02d4;
  localparam int LDPC_ENC_CODEWRD_141_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_141_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_141_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_141_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_141_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_141_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_141_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_141_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_141_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_142_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_142_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_142_BYTE_OFFSET = 13'h02d8;
  localparam int LDPC_ENC_CODEWRD_142_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_142_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_142_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_142_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_142_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_142_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_142_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_142_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_142_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_143_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_143_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_143_BYTE_OFFSET = 13'h02dc;
  localparam int LDPC_ENC_CODEWRD_143_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_143_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_143_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_143_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_143_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_143_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_143_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_143_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_143_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_144_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_144_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_144_BYTE_OFFSET = 13'h02e0;
  localparam int LDPC_ENC_CODEWRD_144_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_144_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_144_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_144_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_144_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_144_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_144_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_144_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_144_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_145_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_145_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_145_BYTE_OFFSET = 13'h02e4;
  localparam int LDPC_ENC_CODEWRD_145_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_145_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_145_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_145_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_145_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_145_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_145_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_145_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_145_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_146_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_146_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_146_BYTE_OFFSET = 13'h02e8;
  localparam int LDPC_ENC_CODEWRD_146_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_146_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_146_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_146_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_146_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_146_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_146_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_146_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_146_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_147_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_147_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_147_BYTE_OFFSET = 13'h02ec;
  localparam int LDPC_ENC_CODEWRD_147_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_147_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_147_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_147_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_147_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_147_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_147_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_147_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_147_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_148_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_148_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_148_BYTE_OFFSET = 13'h02f0;
  localparam int LDPC_ENC_CODEWRD_148_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_148_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_148_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_148_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_148_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_148_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_148_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_148_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_148_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_149_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_149_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_149_BYTE_OFFSET = 13'h02f4;
  localparam int LDPC_ENC_CODEWRD_149_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_149_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_149_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_149_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_149_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_149_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_149_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_149_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_149_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_150_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_150_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_150_BYTE_OFFSET = 13'h02f8;
  localparam int LDPC_ENC_CODEWRD_150_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_150_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_150_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_150_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_150_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_150_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_150_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_150_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_150_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_151_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_151_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_151_BYTE_OFFSET = 13'h02fc;
  localparam int LDPC_ENC_CODEWRD_151_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_151_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_151_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_151_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_151_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_151_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_151_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_151_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_151_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_152_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_152_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_152_BYTE_OFFSET = 13'h0300;
  localparam int LDPC_ENC_CODEWRD_152_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_152_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_152_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_152_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_152_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_152_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_152_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_152_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_152_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_153_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_153_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_153_BYTE_OFFSET = 13'h0304;
  localparam int LDPC_ENC_CODEWRD_153_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_153_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_153_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_153_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_153_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_153_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_153_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_153_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_153_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_154_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_154_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_154_BYTE_OFFSET = 13'h0308;
  localparam int LDPC_ENC_CODEWRD_154_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_154_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_154_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_154_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_154_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_154_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_154_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_154_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_154_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_155_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_155_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_155_BYTE_OFFSET = 13'h030c;
  localparam int LDPC_ENC_CODEWRD_155_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_155_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_155_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_155_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_155_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_155_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_155_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_155_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_155_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_156_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_156_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_156_BYTE_OFFSET = 13'h0310;
  localparam int LDPC_ENC_CODEWRD_156_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_156_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_156_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_156_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_156_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_156_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_156_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_156_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_156_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_157_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_157_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_157_BYTE_OFFSET = 13'h0314;
  localparam int LDPC_ENC_CODEWRD_157_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_157_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_157_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_157_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_157_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_157_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_157_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_157_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_157_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_158_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_158_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_158_BYTE_OFFSET = 13'h0318;
  localparam int LDPC_ENC_CODEWRD_158_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_158_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_158_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_158_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_158_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_158_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_158_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_158_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_158_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_159_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_159_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_159_BYTE_OFFSET = 13'h031c;
  localparam int LDPC_ENC_CODEWRD_159_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_159_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_159_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_159_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_159_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_159_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_159_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_159_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_159_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_160_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_160_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_160_BYTE_OFFSET = 13'h0320;
  localparam int LDPC_ENC_CODEWRD_160_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_160_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_160_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_160_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_160_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_160_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_160_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_160_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_160_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_161_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_161_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_161_BYTE_OFFSET = 13'h0324;
  localparam int LDPC_ENC_CODEWRD_161_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_161_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_161_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_161_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_161_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_161_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_161_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_161_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_161_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_162_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_162_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_162_BYTE_OFFSET = 13'h0328;
  localparam int LDPC_ENC_CODEWRD_162_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_162_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_162_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_162_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_162_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_162_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_162_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_162_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_162_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_163_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_163_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_163_BYTE_OFFSET = 13'h032c;
  localparam int LDPC_ENC_CODEWRD_163_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_163_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_163_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_163_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_163_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_163_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_163_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_163_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_163_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_164_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_164_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_164_BYTE_OFFSET = 13'h0330;
  localparam int LDPC_ENC_CODEWRD_164_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_164_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_164_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_164_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_164_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_164_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_164_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_164_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_164_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_165_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_165_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_165_BYTE_OFFSET = 13'h0334;
  localparam int LDPC_ENC_CODEWRD_165_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_165_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_165_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_165_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_165_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_165_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_165_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_165_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_165_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_166_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_166_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_166_BYTE_OFFSET = 13'h0338;
  localparam int LDPC_ENC_CODEWRD_166_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_166_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_166_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_166_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_166_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_166_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_166_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_166_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_166_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_167_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_167_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_167_BYTE_OFFSET = 13'h033c;
  localparam int LDPC_ENC_CODEWRD_167_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_167_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_167_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_167_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_167_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_167_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_167_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_167_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_167_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_168_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_168_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_168_BYTE_OFFSET = 13'h0340;
  localparam int LDPC_ENC_CODEWRD_168_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_168_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_168_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_168_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_168_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_168_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_168_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_168_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_168_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_169_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_169_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_169_BYTE_OFFSET = 13'h0344;
  localparam int LDPC_ENC_CODEWRD_169_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_169_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_169_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_169_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_169_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_169_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_169_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_169_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_169_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_170_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_170_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_170_BYTE_OFFSET = 13'h0348;
  localparam int LDPC_ENC_CODEWRD_170_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_170_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_170_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_170_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_170_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_170_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_170_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_170_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_170_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_171_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_171_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_171_BYTE_OFFSET = 13'h034c;
  localparam int LDPC_ENC_CODEWRD_171_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_171_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_171_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_171_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_171_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_171_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_171_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_171_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_171_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_172_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_172_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_172_BYTE_OFFSET = 13'h0350;
  localparam int LDPC_ENC_CODEWRD_172_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_172_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_172_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_172_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_172_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_172_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_172_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_172_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_172_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_173_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_173_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_173_BYTE_OFFSET = 13'h0354;
  localparam int LDPC_ENC_CODEWRD_173_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_173_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_173_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_173_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_173_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_173_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_173_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_173_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_173_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_174_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_174_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_174_BYTE_OFFSET = 13'h0358;
  localparam int LDPC_ENC_CODEWRD_174_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_174_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_174_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_174_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_174_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_174_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_174_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_174_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_174_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_175_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_175_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_175_BYTE_OFFSET = 13'h035c;
  localparam int LDPC_ENC_CODEWRD_175_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_175_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_175_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_175_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_175_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_175_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_175_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_175_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_175_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_176_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_176_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_176_BYTE_OFFSET = 13'h0360;
  localparam int LDPC_ENC_CODEWRD_176_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_176_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_176_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_176_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_176_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_176_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_176_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_176_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_176_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_177_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_177_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_177_BYTE_OFFSET = 13'h0364;
  localparam int LDPC_ENC_CODEWRD_177_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_177_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_177_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_177_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_177_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_177_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_177_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_177_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_177_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_178_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_178_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_178_BYTE_OFFSET = 13'h0368;
  localparam int LDPC_ENC_CODEWRD_178_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_178_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_178_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_178_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_178_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_178_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_178_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_178_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_178_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_179_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_179_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_179_BYTE_OFFSET = 13'h036c;
  localparam int LDPC_ENC_CODEWRD_179_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_179_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_179_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_179_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_179_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_179_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_179_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_179_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_179_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_180_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_180_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_180_BYTE_OFFSET = 13'h0370;
  localparam int LDPC_ENC_CODEWRD_180_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_180_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_180_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_180_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_180_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_180_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_180_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_180_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_180_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_181_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_181_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_181_BYTE_OFFSET = 13'h0374;
  localparam int LDPC_ENC_CODEWRD_181_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_181_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_181_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_181_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_181_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_181_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_181_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_181_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_181_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_182_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_182_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_182_BYTE_OFFSET = 13'h0378;
  localparam int LDPC_ENC_CODEWRD_182_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_182_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_182_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_182_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_182_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_182_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_182_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_182_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_182_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_183_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_183_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_183_BYTE_OFFSET = 13'h037c;
  localparam int LDPC_ENC_CODEWRD_183_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_183_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_183_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_183_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_183_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_183_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_183_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_183_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_183_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_184_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_184_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_184_BYTE_OFFSET = 13'h0380;
  localparam int LDPC_ENC_CODEWRD_184_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_184_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_184_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_184_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_184_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_184_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_184_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_184_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_184_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_185_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_185_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_185_BYTE_OFFSET = 13'h0384;
  localparam int LDPC_ENC_CODEWRD_185_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_185_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_185_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_185_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_185_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_185_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_185_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_185_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_185_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_186_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_186_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_186_BYTE_OFFSET = 13'h0388;
  localparam int LDPC_ENC_CODEWRD_186_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_186_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_186_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_186_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_186_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_186_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_186_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_186_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_186_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_187_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_187_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_187_BYTE_OFFSET = 13'h038c;
  localparam int LDPC_ENC_CODEWRD_187_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_187_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_187_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_187_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_187_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_187_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_187_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_187_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_187_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_188_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_188_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_188_BYTE_OFFSET = 13'h0390;
  localparam int LDPC_ENC_CODEWRD_188_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_188_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_188_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_188_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_188_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_188_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_188_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_188_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_188_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_189_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_189_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_189_BYTE_OFFSET = 13'h0394;
  localparam int LDPC_ENC_CODEWRD_189_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_189_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_189_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_189_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_189_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_189_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_189_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_189_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_189_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_190_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_190_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_190_BYTE_OFFSET = 13'h0398;
  localparam int LDPC_ENC_CODEWRD_190_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_190_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_190_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_190_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_190_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_190_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_190_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_190_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_190_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_191_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_191_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_191_BYTE_OFFSET = 13'h039c;
  localparam int LDPC_ENC_CODEWRD_191_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_191_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_191_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_191_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_191_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_191_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_191_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_191_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_191_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_192_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_192_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_192_BYTE_OFFSET = 13'h03a0;
  localparam int LDPC_ENC_CODEWRD_192_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_192_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_192_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_192_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_192_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_192_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_192_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_192_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_192_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_193_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_193_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_193_BYTE_OFFSET = 13'h03a4;
  localparam int LDPC_ENC_CODEWRD_193_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_193_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_193_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_193_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_193_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_193_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_193_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_193_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_193_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_194_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_194_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_194_BYTE_OFFSET = 13'h03a8;
  localparam int LDPC_ENC_CODEWRD_194_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_194_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_194_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_194_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_194_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_194_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_194_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_194_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_194_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_195_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_195_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_195_BYTE_OFFSET = 13'h03ac;
  localparam int LDPC_ENC_CODEWRD_195_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_195_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_195_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_195_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_195_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_195_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_195_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_195_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_195_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_196_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_196_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_196_BYTE_OFFSET = 13'h03b0;
  localparam int LDPC_ENC_CODEWRD_196_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_196_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_196_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_196_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_196_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_196_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_196_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_196_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_196_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_197_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_197_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_197_BYTE_OFFSET = 13'h03b4;
  localparam int LDPC_ENC_CODEWRD_197_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_197_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_197_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_197_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_197_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_197_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_197_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_197_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_197_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_198_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_198_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_198_BYTE_OFFSET = 13'h03b8;
  localparam int LDPC_ENC_CODEWRD_198_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_198_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_198_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_198_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_198_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_198_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_198_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_198_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_198_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_199_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_199_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_199_BYTE_OFFSET = 13'h03bc;
  localparam int LDPC_ENC_CODEWRD_199_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_199_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_199_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_199_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_199_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_199_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_199_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_199_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_199_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_200_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_200_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_200_BYTE_OFFSET = 13'h03c0;
  localparam int LDPC_ENC_CODEWRD_200_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_200_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_200_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_200_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_200_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_200_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_200_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_200_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_200_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_201_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_201_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_201_BYTE_OFFSET = 13'h03c4;
  localparam int LDPC_ENC_CODEWRD_201_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_201_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_201_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_201_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_201_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_201_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_201_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_201_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_201_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_202_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_202_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_202_BYTE_OFFSET = 13'h03c8;
  localparam int LDPC_ENC_CODEWRD_202_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_202_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_202_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_202_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_202_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_202_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_202_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_202_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_202_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_203_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_203_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_203_BYTE_OFFSET = 13'h03cc;
  localparam int LDPC_ENC_CODEWRD_203_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_203_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_203_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_203_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_203_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_203_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_203_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_203_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_203_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_204_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_204_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_204_BYTE_OFFSET = 13'h03d0;
  localparam int LDPC_ENC_CODEWRD_204_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_204_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_204_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_204_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_204_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_204_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_204_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_204_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_204_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_205_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_205_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_205_BYTE_OFFSET = 13'h03d4;
  localparam int LDPC_ENC_CODEWRD_205_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_205_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_205_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_205_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_205_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_205_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_205_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_205_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_205_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_206_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_206_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_206_BYTE_OFFSET = 13'h03d8;
  localparam int LDPC_ENC_CODEWRD_206_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_206_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_206_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_206_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_206_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_206_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_206_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_206_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_206_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_207_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_207_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_207_BYTE_OFFSET = 13'h03dc;
  localparam int LDPC_ENC_CODEWRD_207_ENC_CODEWRDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_207_ENC_CODEWRDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_207_ENC_CODEWRDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_207_ENC_CODEWRDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_207_ENC_CODEWRDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_207_ENC_CODEWRDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_207_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_207_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_207_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_ENC_CODEWRD_VLD_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_VLD_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_VLD_BYTE_OFFSET = 13'h03e0;
  localparam int LDPC_ENC_CODEWRD_VLD_ENC_VALID_CWORDR_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_VLD_ENC_VALID_CWORDR_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_VLD_ENC_VALID_CWORDR_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_VLD_ENC_VALID_CWORDW_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_VLD_ENC_VALID_CWORDW_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_VLD_ENC_VALID_CWORDW_BIT_OFFSET = 1;
  localparam int LDPC_ENC_CODEWRD_VLD_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_ENC_CODEWRD_VLD_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_ENC_CODEWRD_VLD_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_0_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_0_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_0_BYTE_OFFSET = 13'h03e4;
  localparam int LDPC_DEC_CODEWRD_0_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_0_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_0_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_0_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_0_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_0_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_0_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_0_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_0_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_1_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_1_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_1_BYTE_OFFSET = 13'h03e8;
  localparam int LDPC_DEC_CODEWRD_1_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_1_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_1_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_1_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_1_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_1_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_1_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_1_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_1_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_2_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_2_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_2_BYTE_OFFSET = 13'h03ec;
  localparam int LDPC_DEC_CODEWRD_2_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_2_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_2_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_2_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_2_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_2_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_2_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_2_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_2_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_3_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_3_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_3_BYTE_OFFSET = 13'h03f0;
  localparam int LDPC_DEC_CODEWRD_3_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_3_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_3_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_3_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_3_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_3_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_3_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_3_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_3_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_4_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_4_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_4_BYTE_OFFSET = 13'h03f4;
  localparam int LDPC_DEC_CODEWRD_4_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_4_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_4_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_4_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_4_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_4_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_4_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_4_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_4_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_5_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_5_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_5_BYTE_OFFSET = 13'h03f8;
  localparam int LDPC_DEC_CODEWRD_5_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_5_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_5_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_5_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_5_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_5_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_5_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_5_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_5_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_6_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_6_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_6_BYTE_OFFSET = 13'h03fc;
  localparam int LDPC_DEC_CODEWRD_6_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_6_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_6_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_6_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_6_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_6_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_6_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_6_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_6_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_7_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_7_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_7_BYTE_OFFSET = 13'h0400;
  localparam int LDPC_DEC_CODEWRD_7_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_7_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_7_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_7_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_7_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_7_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_7_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_7_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_7_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_8_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_8_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_8_BYTE_OFFSET = 13'h0404;
  localparam int LDPC_DEC_CODEWRD_8_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_8_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_8_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_8_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_8_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_8_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_8_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_8_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_8_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_9_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_9_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_9_BYTE_OFFSET = 13'h0408;
  localparam int LDPC_DEC_CODEWRD_9_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_9_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_9_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_9_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_9_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_9_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_9_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_9_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_9_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_10_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_10_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_10_BYTE_OFFSET = 13'h040c;
  localparam int LDPC_DEC_CODEWRD_10_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_10_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_10_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_10_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_10_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_10_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_10_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_10_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_10_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_11_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_11_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_11_BYTE_OFFSET = 13'h0410;
  localparam int LDPC_DEC_CODEWRD_11_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_11_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_11_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_11_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_11_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_11_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_11_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_11_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_11_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_12_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_12_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_12_BYTE_OFFSET = 13'h0414;
  localparam int LDPC_DEC_CODEWRD_12_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_12_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_12_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_12_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_12_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_12_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_12_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_12_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_12_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_13_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_13_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_13_BYTE_OFFSET = 13'h0418;
  localparam int LDPC_DEC_CODEWRD_13_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_13_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_13_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_13_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_13_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_13_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_13_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_13_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_13_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_14_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_14_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_14_BYTE_OFFSET = 13'h041c;
  localparam int LDPC_DEC_CODEWRD_14_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_14_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_14_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_14_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_14_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_14_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_14_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_14_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_14_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_15_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_15_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_15_BYTE_OFFSET = 13'h0420;
  localparam int LDPC_DEC_CODEWRD_15_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_15_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_15_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_15_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_15_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_15_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_15_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_15_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_15_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_16_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_16_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_16_BYTE_OFFSET = 13'h0424;
  localparam int LDPC_DEC_CODEWRD_16_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_16_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_16_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_16_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_16_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_16_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_16_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_16_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_16_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_17_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_17_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_17_BYTE_OFFSET = 13'h0428;
  localparam int LDPC_DEC_CODEWRD_17_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_17_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_17_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_17_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_17_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_17_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_17_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_17_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_17_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_18_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_18_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_18_BYTE_OFFSET = 13'h042c;
  localparam int LDPC_DEC_CODEWRD_18_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_18_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_18_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_18_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_18_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_18_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_18_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_18_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_18_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_19_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_19_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_19_BYTE_OFFSET = 13'h0430;
  localparam int LDPC_DEC_CODEWRD_19_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_19_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_19_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_19_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_19_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_19_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_19_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_19_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_19_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_20_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_20_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_20_BYTE_OFFSET = 13'h0434;
  localparam int LDPC_DEC_CODEWRD_20_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_20_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_20_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_20_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_20_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_20_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_20_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_20_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_20_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_21_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_21_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_21_BYTE_OFFSET = 13'h0438;
  localparam int LDPC_DEC_CODEWRD_21_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_21_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_21_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_21_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_21_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_21_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_21_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_21_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_21_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_22_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_22_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_22_BYTE_OFFSET = 13'h043c;
  localparam int LDPC_DEC_CODEWRD_22_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_22_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_22_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_22_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_22_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_22_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_22_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_22_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_22_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_23_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_23_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_23_BYTE_OFFSET = 13'h0440;
  localparam int LDPC_DEC_CODEWRD_23_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_23_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_23_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_23_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_23_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_23_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_23_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_23_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_23_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_24_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_24_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_24_BYTE_OFFSET = 13'h0444;
  localparam int LDPC_DEC_CODEWRD_24_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_24_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_24_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_24_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_24_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_24_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_24_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_24_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_24_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_25_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_25_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_25_BYTE_OFFSET = 13'h0448;
  localparam int LDPC_DEC_CODEWRD_25_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_25_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_25_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_25_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_25_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_25_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_25_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_25_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_25_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_26_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_26_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_26_BYTE_OFFSET = 13'h044c;
  localparam int LDPC_DEC_CODEWRD_26_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_26_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_26_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_26_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_26_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_26_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_26_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_26_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_26_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_27_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_27_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_27_BYTE_OFFSET = 13'h0450;
  localparam int LDPC_DEC_CODEWRD_27_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_27_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_27_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_27_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_27_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_27_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_27_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_27_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_27_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_28_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_28_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_28_BYTE_OFFSET = 13'h0454;
  localparam int LDPC_DEC_CODEWRD_28_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_28_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_28_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_28_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_28_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_28_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_28_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_28_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_28_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_29_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_29_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_29_BYTE_OFFSET = 13'h0458;
  localparam int LDPC_DEC_CODEWRD_29_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_29_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_29_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_29_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_29_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_29_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_29_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_29_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_29_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_30_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_30_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_30_BYTE_OFFSET = 13'h045c;
  localparam int LDPC_DEC_CODEWRD_30_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_30_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_30_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_30_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_30_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_30_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_30_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_30_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_30_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_31_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_31_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_31_BYTE_OFFSET = 13'h0460;
  localparam int LDPC_DEC_CODEWRD_31_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_31_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_31_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_31_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_31_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_31_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_31_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_31_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_31_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_32_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_32_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_32_BYTE_OFFSET = 13'h0464;
  localparam int LDPC_DEC_CODEWRD_32_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_32_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_32_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_32_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_32_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_32_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_32_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_32_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_32_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_33_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_33_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_33_BYTE_OFFSET = 13'h0468;
  localparam int LDPC_DEC_CODEWRD_33_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_33_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_33_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_33_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_33_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_33_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_33_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_33_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_33_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_34_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_34_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_34_BYTE_OFFSET = 13'h046c;
  localparam int LDPC_DEC_CODEWRD_34_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_34_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_34_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_34_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_34_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_34_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_34_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_34_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_34_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_35_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_35_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_35_BYTE_OFFSET = 13'h0470;
  localparam int LDPC_DEC_CODEWRD_35_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_35_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_35_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_35_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_35_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_35_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_35_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_35_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_35_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_36_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_36_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_36_BYTE_OFFSET = 13'h0474;
  localparam int LDPC_DEC_CODEWRD_36_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_36_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_36_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_36_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_36_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_36_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_36_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_36_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_36_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_37_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_37_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_37_BYTE_OFFSET = 13'h0478;
  localparam int LDPC_DEC_CODEWRD_37_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_37_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_37_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_37_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_37_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_37_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_37_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_37_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_37_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_38_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_38_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_38_BYTE_OFFSET = 13'h047c;
  localparam int LDPC_DEC_CODEWRD_38_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_38_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_38_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_38_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_38_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_38_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_38_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_38_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_38_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_39_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_39_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_39_BYTE_OFFSET = 13'h0480;
  localparam int LDPC_DEC_CODEWRD_39_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_39_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_39_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_39_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_39_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_39_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_39_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_39_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_39_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_40_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_40_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_40_BYTE_OFFSET = 13'h0484;
  localparam int LDPC_DEC_CODEWRD_40_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_40_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_40_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_40_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_40_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_40_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_40_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_40_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_40_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_41_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_41_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_41_BYTE_OFFSET = 13'h0488;
  localparam int LDPC_DEC_CODEWRD_41_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_41_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_41_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_41_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_41_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_41_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_41_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_41_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_41_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_42_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_42_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_42_BYTE_OFFSET = 13'h048c;
  localparam int LDPC_DEC_CODEWRD_42_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_42_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_42_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_42_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_42_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_42_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_42_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_42_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_42_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_43_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_43_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_43_BYTE_OFFSET = 13'h0490;
  localparam int LDPC_DEC_CODEWRD_43_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_43_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_43_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_43_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_43_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_43_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_43_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_43_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_43_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_44_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_44_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_44_BYTE_OFFSET = 13'h0494;
  localparam int LDPC_DEC_CODEWRD_44_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_44_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_44_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_44_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_44_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_44_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_44_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_44_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_44_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_45_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_45_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_45_BYTE_OFFSET = 13'h0498;
  localparam int LDPC_DEC_CODEWRD_45_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_45_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_45_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_45_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_45_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_45_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_45_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_45_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_45_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_46_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_46_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_46_BYTE_OFFSET = 13'h049c;
  localparam int LDPC_DEC_CODEWRD_46_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_46_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_46_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_46_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_46_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_46_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_46_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_46_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_46_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_47_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_47_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_47_BYTE_OFFSET = 13'h04a0;
  localparam int LDPC_DEC_CODEWRD_47_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_47_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_47_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_47_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_47_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_47_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_47_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_47_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_47_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_48_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_48_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_48_BYTE_OFFSET = 13'h04a4;
  localparam int LDPC_DEC_CODEWRD_48_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_48_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_48_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_48_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_48_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_48_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_48_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_48_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_48_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_49_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_49_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_49_BYTE_OFFSET = 13'h04a8;
  localparam int LDPC_DEC_CODEWRD_49_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_49_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_49_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_49_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_49_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_49_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_49_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_49_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_49_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_50_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_50_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_50_BYTE_OFFSET = 13'h04ac;
  localparam int LDPC_DEC_CODEWRD_50_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_50_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_50_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_50_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_50_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_50_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_50_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_50_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_50_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_51_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_51_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_51_BYTE_OFFSET = 13'h04b0;
  localparam int LDPC_DEC_CODEWRD_51_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_51_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_51_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_51_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_51_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_51_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_51_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_51_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_51_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_52_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_52_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_52_BYTE_OFFSET = 13'h04b4;
  localparam int LDPC_DEC_CODEWRD_52_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_52_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_52_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_52_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_52_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_52_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_52_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_52_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_52_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_53_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_53_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_53_BYTE_OFFSET = 13'h04b8;
  localparam int LDPC_DEC_CODEWRD_53_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_53_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_53_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_53_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_53_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_53_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_53_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_53_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_53_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_54_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_54_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_54_BYTE_OFFSET = 13'h04bc;
  localparam int LDPC_DEC_CODEWRD_54_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_54_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_54_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_54_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_54_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_54_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_54_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_54_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_54_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_55_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_55_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_55_BYTE_OFFSET = 13'h04c0;
  localparam int LDPC_DEC_CODEWRD_55_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_55_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_55_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_55_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_55_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_55_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_55_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_55_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_55_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_56_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_56_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_56_BYTE_OFFSET = 13'h04c4;
  localparam int LDPC_DEC_CODEWRD_56_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_56_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_56_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_56_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_56_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_56_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_56_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_56_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_56_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_57_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_57_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_57_BYTE_OFFSET = 13'h04c8;
  localparam int LDPC_DEC_CODEWRD_57_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_57_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_57_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_57_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_57_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_57_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_57_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_57_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_57_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_58_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_58_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_58_BYTE_OFFSET = 13'h04cc;
  localparam int LDPC_DEC_CODEWRD_58_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_58_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_58_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_58_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_58_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_58_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_58_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_58_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_58_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_59_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_59_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_59_BYTE_OFFSET = 13'h04d0;
  localparam int LDPC_DEC_CODEWRD_59_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_59_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_59_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_59_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_59_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_59_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_59_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_59_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_59_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_60_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_60_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_60_BYTE_OFFSET = 13'h04d4;
  localparam int LDPC_DEC_CODEWRD_60_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_60_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_60_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_60_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_60_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_60_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_60_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_60_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_60_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_61_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_61_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_61_BYTE_OFFSET = 13'h04d8;
  localparam int LDPC_DEC_CODEWRD_61_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_61_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_61_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_61_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_61_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_61_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_61_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_61_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_61_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_62_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_62_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_62_BYTE_OFFSET = 13'h04dc;
  localparam int LDPC_DEC_CODEWRD_62_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_62_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_62_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_62_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_62_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_62_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_62_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_62_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_62_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_63_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_63_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_63_BYTE_OFFSET = 13'h04e0;
  localparam int LDPC_DEC_CODEWRD_63_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_63_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_63_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_63_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_63_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_63_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_63_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_63_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_63_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_64_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_64_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_64_BYTE_OFFSET = 13'h04e4;
  localparam int LDPC_DEC_CODEWRD_64_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_64_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_64_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_64_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_64_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_64_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_64_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_64_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_64_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_65_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_65_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_65_BYTE_OFFSET = 13'h04e8;
  localparam int LDPC_DEC_CODEWRD_65_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_65_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_65_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_65_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_65_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_65_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_65_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_65_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_65_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_66_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_66_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_66_BYTE_OFFSET = 13'h04ec;
  localparam int LDPC_DEC_CODEWRD_66_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_66_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_66_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_66_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_66_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_66_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_66_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_66_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_66_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_67_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_67_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_67_BYTE_OFFSET = 13'h04f0;
  localparam int LDPC_DEC_CODEWRD_67_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_67_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_67_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_67_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_67_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_67_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_67_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_67_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_67_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_68_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_68_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_68_BYTE_OFFSET = 13'h04f4;
  localparam int LDPC_DEC_CODEWRD_68_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_68_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_68_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_68_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_68_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_68_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_68_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_68_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_68_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_69_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_69_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_69_BYTE_OFFSET = 13'h04f8;
  localparam int LDPC_DEC_CODEWRD_69_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_69_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_69_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_69_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_69_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_69_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_69_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_69_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_69_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_70_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_70_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_70_BYTE_OFFSET = 13'h04fc;
  localparam int LDPC_DEC_CODEWRD_70_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_70_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_70_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_70_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_70_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_70_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_70_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_70_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_70_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_71_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_71_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_71_BYTE_OFFSET = 13'h0500;
  localparam int LDPC_DEC_CODEWRD_71_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_71_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_71_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_71_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_71_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_71_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_71_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_71_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_71_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_72_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_72_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_72_BYTE_OFFSET = 13'h0504;
  localparam int LDPC_DEC_CODEWRD_72_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_72_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_72_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_72_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_72_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_72_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_72_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_72_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_72_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_73_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_73_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_73_BYTE_OFFSET = 13'h0508;
  localparam int LDPC_DEC_CODEWRD_73_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_73_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_73_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_73_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_73_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_73_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_73_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_73_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_73_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_74_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_74_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_74_BYTE_OFFSET = 13'h050c;
  localparam int LDPC_DEC_CODEWRD_74_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_74_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_74_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_74_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_74_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_74_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_74_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_74_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_74_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_75_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_75_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_75_BYTE_OFFSET = 13'h0510;
  localparam int LDPC_DEC_CODEWRD_75_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_75_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_75_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_75_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_75_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_75_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_75_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_75_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_75_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_76_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_76_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_76_BYTE_OFFSET = 13'h0514;
  localparam int LDPC_DEC_CODEWRD_76_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_76_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_76_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_76_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_76_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_76_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_76_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_76_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_76_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_77_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_77_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_77_BYTE_OFFSET = 13'h0518;
  localparam int LDPC_DEC_CODEWRD_77_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_77_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_77_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_77_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_77_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_77_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_77_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_77_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_77_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_78_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_78_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_78_BYTE_OFFSET = 13'h051c;
  localparam int LDPC_DEC_CODEWRD_78_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_78_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_78_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_78_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_78_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_78_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_78_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_78_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_78_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_79_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_79_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_79_BYTE_OFFSET = 13'h0520;
  localparam int LDPC_DEC_CODEWRD_79_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_79_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_79_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_79_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_79_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_79_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_79_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_79_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_79_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_80_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_80_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_80_BYTE_OFFSET = 13'h0524;
  localparam int LDPC_DEC_CODEWRD_80_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_80_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_80_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_80_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_80_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_80_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_80_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_80_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_80_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_81_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_81_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_81_BYTE_OFFSET = 13'h0528;
  localparam int LDPC_DEC_CODEWRD_81_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_81_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_81_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_81_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_81_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_81_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_81_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_81_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_81_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_82_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_82_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_82_BYTE_OFFSET = 13'h052c;
  localparam int LDPC_DEC_CODEWRD_82_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_82_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_82_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_82_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_82_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_82_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_82_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_82_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_82_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_83_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_83_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_83_BYTE_OFFSET = 13'h0530;
  localparam int LDPC_DEC_CODEWRD_83_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_83_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_83_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_83_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_83_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_83_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_83_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_83_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_83_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_84_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_84_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_84_BYTE_OFFSET = 13'h0534;
  localparam int LDPC_DEC_CODEWRD_84_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_84_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_84_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_84_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_84_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_84_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_84_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_84_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_84_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_85_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_85_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_85_BYTE_OFFSET = 13'h0538;
  localparam int LDPC_DEC_CODEWRD_85_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_85_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_85_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_85_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_85_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_85_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_85_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_85_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_85_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_86_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_86_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_86_BYTE_OFFSET = 13'h053c;
  localparam int LDPC_DEC_CODEWRD_86_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_86_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_86_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_86_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_86_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_86_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_86_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_86_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_86_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_87_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_87_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_87_BYTE_OFFSET = 13'h0540;
  localparam int LDPC_DEC_CODEWRD_87_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_87_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_87_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_87_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_87_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_87_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_87_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_87_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_87_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_88_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_88_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_88_BYTE_OFFSET = 13'h0544;
  localparam int LDPC_DEC_CODEWRD_88_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_88_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_88_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_88_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_88_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_88_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_88_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_88_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_88_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_89_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_89_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_89_BYTE_OFFSET = 13'h0548;
  localparam int LDPC_DEC_CODEWRD_89_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_89_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_89_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_89_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_89_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_89_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_89_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_89_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_89_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_90_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_90_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_90_BYTE_OFFSET = 13'h054c;
  localparam int LDPC_DEC_CODEWRD_90_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_90_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_90_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_90_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_90_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_90_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_90_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_90_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_90_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_91_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_91_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_91_BYTE_OFFSET = 13'h0550;
  localparam int LDPC_DEC_CODEWRD_91_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_91_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_91_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_91_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_91_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_91_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_91_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_91_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_91_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_92_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_92_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_92_BYTE_OFFSET = 13'h0554;
  localparam int LDPC_DEC_CODEWRD_92_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_92_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_92_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_92_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_92_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_92_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_92_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_92_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_92_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_93_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_93_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_93_BYTE_OFFSET = 13'h0558;
  localparam int LDPC_DEC_CODEWRD_93_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_93_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_93_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_93_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_93_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_93_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_93_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_93_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_93_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_94_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_94_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_94_BYTE_OFFSET = 13'h055c;
  localparam int LDPC_DEC_CODEWRD_94_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_94_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_94_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_94_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_94_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_94_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_94_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_94_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_94_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_95_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_95_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_95_BYTE_OFFSET = 13'h0560;
  localparam int LDPC_DEC_CODEWRD_95_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_95_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_95_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_95_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_95_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_95_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_95_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_95_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_95_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_96_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_96_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_96_BYTE_OFFSET = 13'h0564;
  localparam int LDPC_DEC_CODEWRD_96_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_96_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_96_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_96_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_96_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_96_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_96_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_96_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_96_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_97_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_97_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_97_BYTE_OFFSET = 13'h0568;
  localparam int LDPC_DEC_CODEWRD_97_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_97_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_97_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_97_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_97_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_97_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_97_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_97_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_97_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_98_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_98_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_98_BYTE_OFFSET = 13'h056c;
  localparam int LDPC_DEC_CODEWRD_98_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_98_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_98_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_98_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_98_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_98_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_98_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_98_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_98_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_99_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_99_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_99_BYTE_OFFSET = 13'h0570;
  localparam int LDPC_DEC_CODEWRD_99_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_99_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_99_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_99_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_99_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_99_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_99_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_99_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_99_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_100_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_100_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_100_BYTE_OFFSET = 13'h0574;
  localparam int LDPC_DEC_CODEWRD_100_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_100_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_100_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_100_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_100_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_100_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_100_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_100_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_100_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_101_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_101_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_101_BYTE_OFFSET = 13'h0578;
  localparam int LDPC_DEC_CODEWRD_101_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_101_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_101_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_101_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_101_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_101_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_101_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_101_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_101_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_102_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_102_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_102_BYTE_OFFSET = 13'h057c;
  localparam int LDPC_DEC_CODEWRD_102_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_102_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_102_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_102_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_102_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_102_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_102_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_102_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_102_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_103_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_103_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_103_BYTE_OFFSET = 13'h0580;
  localparam int LDPC_DEC_CODEWRD_103_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_103_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_103_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_103_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_103_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_103_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_103_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_103_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_103_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_104_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_104_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_104_BYTE_OFFSET = 13'h0584;
  localparam int LDPC_DEC_CODEWRD_104_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_104_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_104_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_104_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_104_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_104_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_104_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_104_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_104_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_105_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_105_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_105_BYTE_OFFSET = 13'h0588;
  localparam int LDPC_DEC_CODEWRD_105_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_105_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_105_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_105_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_105_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_105_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_105_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_105_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_105_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_106_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_106_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_106_BYTE_OFFSET = 13'h058c;
  localparam int LDPC_DEC_CODEWRD_106_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_106_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_106_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_106_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_106_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_106_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_106_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_106_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_106_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_107_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_107_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_107_BYTE_OFFSET = 13'h0590;
  localparam int LDPC_DEC_CODEWRD_107_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_107_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_107_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_107_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_107_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_107_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_107_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_107_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_107_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_108_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_108_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_108_BYTE_OFFSET = 13'h0594;
  localparam int LDPC_DEC_CODEWRD_108_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_108_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_108_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_108_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_108_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_108_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_108_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_108_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_108_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_109_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_109_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_109_BYTE_OFFSET = 13'h0598;
  localparam int LDPC_DEC_CODEWRD_109_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_109_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_109_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_109_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_109_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_109_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_109_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_109_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_109_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_110_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_110_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_110_BYTE_OFFSET = 13'h059c;
  localparam int LDPC_DEC_CODEWRD_110_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_110_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_110_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_110_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_110_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_110_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_110_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_110_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_110_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_111_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_111_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_111_BYTE_OFFSET = 13'h05a0;
  localparam int LDPC_DEC_CODEWRD_111_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_111_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_111_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_111_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_111_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_111_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_111_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_111_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_111_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_112_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_112_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_112_BYTE_OFFSET = 13'h05a4;
  localparam int LDPC_DEC_CODEWRD_112_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_112_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_112_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_112_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_112_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_112_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_112_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_112_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_112_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_113_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_113_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_113_BYTE_OFFSET = 13'h05a8;
  localparam int LDPC_DEC_CODEWRD_113_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_113_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_113_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_113_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_113_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_113_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_113_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_113_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_113_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_114_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_114_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_114_BYTE_OFFSET = 13'h05ac;
  localparam int LDPC_DEC_CODEWRD_114_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_114_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_114_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_114_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_114_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_114_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_114_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_114_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_114_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_115_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_115_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_115_BYTE_OFFSET = 13'h05b0;
  localparam int LDPC_DEC_CODEWRD_115_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_115_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_115_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_115_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_115_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_115_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_115_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_115_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_115_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_116_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_116_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_116_BYTE_OFFSET = 13'h05b4;
  localparam int LDPC_DEC_CODEWRD_116_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_116_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_116_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_116_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_116_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_116_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_116_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_116_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_116_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_117_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_117_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_117_BYTE_OFFSET = 13'h05b8;
  localparam int LDPC_DEC_CODEWRD_117_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_117_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_117_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_117_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_117_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_117_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_117_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_117_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_117_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_118_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_118_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_118_BYTE_OFFSET = 13'h05bc;
  localparam int LDPC_DEC_CODEWRD_118_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_118_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_118_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_118_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_118_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_118_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_118_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_118_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_118_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_119_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_119_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_119_BYTE_OFFSET = 13'h05c0;
  localparam int LDPC_DEC_CODEWRD_119_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_119_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_119_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_119_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_119_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_119_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_119_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_119_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_119_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_120_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_120_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_120_BYTE_OFFSET = 13'h05c4;
  localparam int LDPC_DEC_CODEWRD_120_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_120_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_120_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_120_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_120_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_120_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_120_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_120_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_120_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_121_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_121_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_121_BYTE_OFFSET = 13'h05c8;
  localparam int LDPC_DEC_CODEWRD_121_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_121_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_121_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_121_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_121_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_121_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_121_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_121_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_121_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_122_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_122_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_122_BYTE_OFFSET = 13'h05cc;
  localparam int LDPC_DEC_CODEWRD_122_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_122_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_122_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_122_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_122_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_122_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_122_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_122_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_122_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_123_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_123_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_123_BYTE_OFFSET = 13'h05d0;
  localparam int LDPC_DEC_CODEWRD_123_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_123_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_123_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_123_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_123_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_123_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_123_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_123_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_123_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_124_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_124_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_124_BYTE_OFFSET = 13'h05d4;
  localparam int LDPC_DEC_CODEWRD_124_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_124_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_124_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_124_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_124_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_124_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_124_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_124_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_124_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_125_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_125_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_125_BYTE_OFFSET = 13'h05d8;
  localparam int LDPC_DEC_CODEWRD_125_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_125_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_125_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_125_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_125_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_125_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_125_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_125_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_125_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_126_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_126_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_126_BYTE_OFFSET = 13'h05dc;
  localparam int LDPC_DEC_CODEWRD_126_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_126_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_126_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_126_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_126_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_126_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_126_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_126_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_126_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_127_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_127_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_127_BYTE_OFFSET = 13'h05e0;
  localparam int LDPC_DEC_CODEWRD_127_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_127_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_127_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_127_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_127_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_127_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_127_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_127_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_127_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_128_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_128_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_128_BYTE_OFFSET = 13'h05e4;
  localparam int LDPC_DEC_CODEWRD_128_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_128_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_128_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_128_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_128_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_128_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_128_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_128_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_128_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_129_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_129_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_129_BYTE_OFFSET = 13'h05e8;
  localparam int LDPC_DEC_CODEWRD_129_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_129_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_129_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_129_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_129_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_129_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_129_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_129_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_129_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_130_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_130_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_130_BYTE_OFFSET = 13'h05ec;
  localparam int LDPC_DEC_CODEWRD_130_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_130_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_130_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_130_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_130_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_130_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_130_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_130_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_130_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_131_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_131_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_131_BYTE_OFFSET = 13'h05f0;
  localparam int LDPC_DEC_CODEWRD_131_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_131_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_131_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_131_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_131_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_131_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_131_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_131_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_131_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_132_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_132_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_132_BYTE_OFFSET = 13'h05f4;
  localparam int LDPC_DEC_CODEWRD_132_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_132_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_132_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_132_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_132_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_132_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_132_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_132_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_132_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_133_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_133_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_133_BYTE_OFFSET = 13'h05f8;
  localparam int LDPC_DEC_CODEWRD_133_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_133_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_133_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_133_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_133_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_133_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_133_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_133_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_133_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_134_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_134_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_134_BYTE_OFFSET = 13'h05fc;
  localparam int LDPC_DEC_CODEWRD_134_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_134_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_134_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_134_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_134_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_134_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_134_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_134_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_134_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_135_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_135_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_135_BYTE_OFFSET = 13'h0600;
  localparam int LDPC_DEC_CODEWRD_135_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_135_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_135_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_135_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_135_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_135_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_135_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_135_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_135_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_136_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_136_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_136_BYTE_OFFSET = 13'h0604;
  localparam int LDPC_DEC_CODEWRD_136_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_136_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_136_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_136_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_136_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_136_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_136_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_136_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_136_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_137_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_137_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_137_BYTE_OFFSET = 13'h0608;
  localparam int LDPC_DEC_CODEWRD_137_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_137_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_137_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_137_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_137_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_137_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_137_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_137_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_137_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_138_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_138_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_138_BYTE_OFFSET = 13'h060c;
  localparam int LDPC_DEC_CODEWRD_138_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_138_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_138_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_138_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_138_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_138_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_138_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_138_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_138_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_139_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_139_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_139_BYTE_OFFSET = 13'h0610;
  localparam int LDPC_DEC_CODEWRD_139_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_139_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_139_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_139_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_139_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_139_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_139_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_139_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_139_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_140_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_140_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_140_BYTE_OFFSET = 13'h0614;
  localparam int LDPC_DEC_CODEWRD_140_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_140_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_140_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_140_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_140_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_140_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_140_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_140_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_140_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_141_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_141_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_141_BYTE_OFFSET = 13'h0618;
  localparam int LDPC_DEC_CODEWRD_141_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_141_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_141_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_141_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_141_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_141_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_141_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_141_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_141_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_142_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_142_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_142_BYTE_OFFSET = 13'h061c;
  localparam int LDPC_DEC_CODEWRD_142_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_142_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_142_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_142_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_142_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_142_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_142_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_142_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_142_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_143_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_143_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_143_BYTE_OFFSET = 13'h0620;
  localparam int LDPC_DEC_CODEWRD_143_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_143_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_143_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_143_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_143_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_143_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_143_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_143_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_143_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_144_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_144_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_144_BYTE_OFFSET = 13'h0624;
  localparam int LDPC_DEC_CODEWRD_144_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_144_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_144_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_144_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_144_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_144_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_144_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_144_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_144_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_145_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_145_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_145_BYTE_OFFSET = 13'h0628;
  localparam int LDPC_DEC_CODEWRD_145_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_145_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_145_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_145_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_145_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_145_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_145_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_145_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_145_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_146_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_146_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_146_BYTE_OFFSET = 13'h062c;
  localparam int LDPC_DEC_CODEWRD_146_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_146_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_146_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_146_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_146_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_146_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_146_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_146_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_146_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_147_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_147_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_147_BYTE_OFFSET = 13'h0630;
  localparam int LDPC_DEC_CODEWRD_147_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_147_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_147_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_147_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_147_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_147_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_147_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_147_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_147_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_148_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_148_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_148_BYTE_OFFSET = 13'h0634;
  localparam int LDPC_DEC_CODEWRD_148_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_148_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_148_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_148_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_148_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_148_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_148_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_148_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_148_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_149_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_149_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_149_BYTE_OFFSET = 13'h0638;
  localparam int LDPC_DEC_CODEWRD_149_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_149_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_149_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_149_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_149_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_149_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_149_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_149_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_149_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_150_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_150_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_150_BYTE_OFFSET = 13'h063c;
  localparam int LDPC_DEC_CODEWRD_150_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_150_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_150_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_150_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_150_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_150_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_150_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_150_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_150_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_151_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_151_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_151_BYTE_OFFSET = 13'h0640;
  localparam int LDPC_DEC_CODEWRD_151_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_151_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_151_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_151_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_151_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_151_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_151_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_151_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_151_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_152_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_152_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_152_BYTE_OFFSET = 13'h0644;
  localparam int LDPC_DEC_CODEWRD_152_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_152_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_152_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_152_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_152_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_152_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_152_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_152_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_152_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_153_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_153_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_153_BYTE_OFFSET = 13'h0648;
  localparam int LDPC_DEC_CODEWRD_153_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_153_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_153_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_153_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_153_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_153_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_153_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_153_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_153_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_154_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_154_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_154_BYTE_OFFSET = 13'h064c;
  localparam int LDPC_DEC_CODEWRD_154_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_154_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_154_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_154_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_154_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_154_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_154_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_154_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_154_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_155_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_155_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_155_BYTE_OFFSET = 13'h0650;
  localparam int LDPC_DEC_CODEWRD_155_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_155_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_155_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_155_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_155_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_155_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_155_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_155_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_155_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_156_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_156_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_156_BYTE_OFFSET = 13'h0654;
  localparam int LDPC_DEC_CODEWRD_156_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_156_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_156_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_156_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_156_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_156_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_156_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_156_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_156_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_157_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_157_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_157_BYTE_OFFSET = 13'h0658;
  localparam int LDPC_DEC_CODEWRD_157_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_157_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_157_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_157_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_157_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_157_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_157_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_157_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_157_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_158_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_158_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_158_BYTE_OFFSET = 13'h065c;
  localparam int LDPC_DEC_CODEWRD_158_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_158_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_158_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_158_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_158_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_158_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_158_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_158_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_158_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_159_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_159_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_159_BYTE_OFFSET = 13'h0660;
  localparam int LDPC_DEC_CODEWRD_159_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_159_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_159_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_159_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_159_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_159_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_159_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_159_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_159_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_160_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_160_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_160_BYTE_OFFSET = 13'h0664;
  localparam int LDPC_DEC_CODEWRD_160_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_160_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_160_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_160_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_160_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_160_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_160_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_160_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_160_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_161_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_161_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_161_BYTE_OFFSET = 13'h0668;
  localparam int LDPC_DEC_CODEWRD_161_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_161_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_161_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_161_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_161_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_161_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_161_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_161_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_161_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_162_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_162_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_162_BYTE_OFFSET = 13'h066c;
  localparam int LDPC_DEC_CODEWRD_162_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_162_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_162_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_162_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_162_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_162_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_162_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_162_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_162_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_163_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_163_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_163_BYTE_OFFSET = 13'h0670;
  localparam int LDPC_DEC_CODEWRD_163_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_163_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_163_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_163_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_163_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_163_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_163_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_163_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_163_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_164_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_164_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_164_BYTE_OFFSET = 13'h0674;
  localparam int LDPC_DEC_CODEWRD_164_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_164_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_164_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_164_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_164_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_164_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_164_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_164_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_164_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_165_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_165_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_165_BYTE_OFFSET = 13'h0678;
  localparam int LDPC_DEC_CODEWRD_165_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_165_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_165_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_165_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_165_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_165_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_165_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_165_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_165_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_166_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_166_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_166_BYTE_OFFSET = 13'h067c;
  localparam int LDPC_DEC_CODEWRD_166_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_166_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_166_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_166_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_166_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_166_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_166_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_166_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_166_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_167_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_167_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_167_BYTE_OFFSET = 13'h0680;
  localparam int LDPC_DEC_CODEWRD_167_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_167_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_167_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_167_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_167_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_167_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_167_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_167_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_167_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_168_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_168_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_168_BYTE_OFFSET = 13'h0684;
  localparam int LDPC_DEC_CODEWRD_168_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_168_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_168_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_168_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_168_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_168_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_168_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_168_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_168_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_169_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_169_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_169_BYTE_OFFSET = 13'h0688;
  localparam int LDPC_DEC_CODEWRD_169_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_169_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_169_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_169_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_169_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_169_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_169_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_169_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_169_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_170_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_170_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_170_BYTE_OFFSET = 13'h068c;
  localparam int LDPC_DEC_CODEWRD_170_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_170_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_170_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_170_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_170_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_170_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_170_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_170_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_170_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_171_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_171_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_171_BYTE_OFFSET = 13'h0690;
  localparam int LDPC_DEC_CODEWRD_171_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_171_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_171_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_171_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_171_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_171_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_171_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_171_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_171_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_172_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_172_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_172_BYTE_OFFSET = 13'h0694;
  localparam int LDPC_DEC_CODEWRD_172_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_172_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_172_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_172_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_172_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_172_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_172_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_172_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_172_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_173_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_173_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_173_BYTE_OFFSET = 13'h0698;
  localparam int LDPC_DEC_CODEWRD_173_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_173_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_173_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_173_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_173_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_173_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_173_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_173_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_173_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_174_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_174_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_174_BYTE_OFFSET = 13'h069c;
  localparam int LDPC_DEC_CODEWRD_174_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_174_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_174_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_174_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_174_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_174_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_174_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_174_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_174_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_175_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_175_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_175_BYTE_OFFSET = 13'h06a0;
  localparam int LDPC_DEC_CODEWRD_175_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_175_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_175_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_175_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_175_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_175_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_175_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_175_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_175_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_176_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_176_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_176_BYTE_OFFSET = 13'h06a4;
  localparam int LDPC_DEC_CODEWRD_176_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_176_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_176_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_176_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_176_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_176_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_176_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_176_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_176_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_177_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_177_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_177_BYTE_OFFSET = 13'h06a8;
  localparam int LDPC_DEC_CODEWRD_177_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_177_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_177_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_177_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_177_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_177_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_177_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_177_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_177_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_178_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_178_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_178_BYTE_OFFSET = 13'h06ac;
  localparam int LDPC_DEC_CODEWRD_178_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_178_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_178_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_178_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_178_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_178_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_178_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_178_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_178_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_179_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_179_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_179_BYTE_OFFSET = 13'h06b0;
  localparam int LDPC_DEC_CODEWRD_179_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_179_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_179_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_179_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_179_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_179_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_179_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_179_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_179_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_180_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_180_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_180_BYTE_OFFSET = 13'h06b4;
  localparam int LDPC_DEC_CODEWRD_180_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_180_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_180_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_180_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_180_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_180_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_180_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_180_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_180_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_181_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_181_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_181_BYTE_OFFSET = 13'h06b8;
  localparam int LDPC_DEC_CODEWRD_181_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_181_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_181_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_181_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_181_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_181_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_181_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_181_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_181_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_182_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_182_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_182_BYTE_OFFSET = 13'h06bc;
  localparam int LDPC_DEC_CODEWRD_182_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_182_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_182_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_182_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_182_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_182_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_182_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_182_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_182_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_183_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_183_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_183_BYTE_OFFSET = 13'h06c0;
  localparam int LDPC_DEC_CODEWRD_183_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_183_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_183_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_183_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_183_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_183_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_183_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_183_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_183_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_184_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_184_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_184_BYTE_OFFSET = 13'h06c4;
  localparam int LDPC_DEC_CODEWRD_184_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_184_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_184_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_184_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_184_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_184_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_184_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_184_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_184_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_185_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_185_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_185_BYTE_OFFSET = 13'h06c8;
  localparam int LDPC_DEC_CODEWRD_185_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_185_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_185_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_185_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_185_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_185_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_185_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_185_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_185_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_186_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_186_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_186_BYTE_OFFSET = 13'h06cc;
  localparam int LDPC_DEC_CODEWRD_186_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_186_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_186_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_186_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_186_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_186_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_186_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_186_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_186_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_187_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_187_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_187_BYTE_OFFSET = 13'h06d0;
  localparam int LDPC_DEC_CODEWRD_187_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_187_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_187_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_187_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_187_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_187_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_187_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_187_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_187_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_188_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_188_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_188_BYTE_OFFSET = 13'h06d4;
  localparam int LDPC_DEC_CODEWRD_188_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_188_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_188_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_188_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_188_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_188_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_188_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_188_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_188_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_189_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_189_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_189_BYTE_OFFSET = 13'h06d8;
  localparam int LDPC_DEC_CODEWRD_189_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_189_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_189_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_189_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_189_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_189_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_189_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_189_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_189_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_190_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_190_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_190_BYTE_OFFSET = 13'h06dc;
  localparam int LDPC_DEC_CODEWRD_190_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_190_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_190_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_190_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_190_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_190_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_190_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_190_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_190_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_191_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_191_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_191_BYTE_OFFSET = 13'h06e0;
  localparam int LDPC_DEC_CODEWRD_191_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_191_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_191_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_191_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_191_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_191_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_191_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_191_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_191_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_192_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_192_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_192_BYTE_OFFSET = 13'h06e4;
  localparam int LDPC_DEC_CODEWRD_192_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_192_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_192_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_192_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_192_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_192_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_192_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_192_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_192_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_193_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_193_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_193_BYTE_OFFSET = 13'h06e8;
  localparam int LDPC_DEC_CODEWRD_193_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_193_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_193_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_193_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_193_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_193_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_193_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_193_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_193_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_194_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_194_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_194_BYTE_OFFSET = 13'h06ec;
  localparam int LDPC_DEC_CODEWRD_194_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_194_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_194_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_194_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_194_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_194_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_194_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_194_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_194_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_195_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_195_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_195_BYTE_OFFSET = 13'h06f0;
  localparam int LDPC_DEC_CODEWRD_195_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_195_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_195_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_195_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_195_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_195_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_195_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_195_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_195_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_196_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_196_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_196_BYTE_OFFSET = 13'h06f4;
  localparam int LDPC_DEC_CODEWRD_196_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_196_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_196_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_196_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_196_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_196_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_196_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_196_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_196_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_197_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_197_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_197_BYTE_OFFSET = 13'h06f8;
  localparam int LDPC_DEC_CODEWRD_197_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_197_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_197_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_197_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_197_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_197_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_197_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_197_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_197_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_198_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_198_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_198_BYTE_OFFSET = 13'h06fc;
  localparam int LDPC_DEC_CODEWRD_198_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_198_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_198_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_198_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_198_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_198_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_198_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_198_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_198_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_199_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_199_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_199_BYTE_OFFSET = 13'h0700;
  localparam int LDPC_DEC_CODEWRD_199_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_199_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_199_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_199_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_199_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_199_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_199_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_199_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_199_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_200_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_200_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_200_BYTE_OFFSET = 13'h0704;
  localparam int LDPC_DEC_CODEWRD_200_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_200_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_200_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_200_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_200_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_200_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_200_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_200_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_200_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_201_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_201_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_201_BYTE_OFFSET = 13'h0708;
  localparam int LDPC_DEC_CODEWRD_201_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_201_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_201_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_201_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_201_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_201_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_201_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_201_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_201_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_202_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_202_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_202_BYTE_OFFSET = 13'h070c;
  localparam int LDPC_DEC_CODEWRD_202_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_202_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_202_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_202_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_202_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_202_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_202_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_202_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_202_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_203_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_203_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_203_BYTE_OFFSET = 13'h0710;
  localparam int LDPC_DEC_CODEWRD_203_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_203_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_203_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_203_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_203_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_203_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_203_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_203_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_203_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_204_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_204_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_204_BYTE_OFFSET = 13'h0714;
  localparam int LDPC_DEC_CODEWRD_204_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_204_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_204_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_204_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_204_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_204_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_204_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_204_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_204_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_205_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_205_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_205_BYTE_OFFSET = 13'h0718;
  localparam int LDPC_DEC_CODEWRD_205_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_205_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_205_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_205_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_205_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_205_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_205_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_205_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_205_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_206_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_206_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_206_BYTE_OFFSET = 13'h071c;
  localparam int LDPC_DEC_CODEWRD_206_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_206_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_206_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_206_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_206_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_206_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_206_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_206_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_206_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_CODEWRD_207_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_207_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_207_BYTE_OFFSET = 13'h0720;
  localparam int LDPC_DEC_CODEWRD_207_CWORD_Q0R_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_207_CWORD_Q0R_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_207_CWORD_Q0R_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_207_CWORD_Q0W_BIT_WIDTH = 2;
  localparam bit [1:0] LDPC_DEC_CODEWRD_207_CWORD_Q0W_BIT_MASK = 2'h3;
  localparam int LDPC_DEC_CODEWRD_207_CWORD_Q0W_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CODEWRD_207_RESERVED_BIT_WIDTH = 28;
  localparam bit [27:0] LDPC_DEC_CODEWRD_207_RESERVED_BIT_MASK = 28'hfffffff;
  localparam int LDPC_DEC_CODEWRD_207_RESERVED_BIT_OFFSET = 4;
  localparam int LDPC_DEC_EXPSYND_0_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_0_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_0_BYTE_OFFSET = 13'h0724;
  localparam int LDPC_DEC_EXPSYND_0_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_0_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_0_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_0_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_0_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_0_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_0_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_0_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_0_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_1_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_1_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_1_BYTE_OFFSET = 13'h0728;
  localparam int LDPC_DEC_EXPSYND_1_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_1_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_1_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_1_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_1_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_1_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_1_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_1_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_1_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_2_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_2_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_2_BYTE_OFFSET = 13'h072c;
  localparam int LDPC_DEC_EXPSYND_2_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_2_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_2_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_2_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_2_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_2_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_2_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_2_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_2_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_3_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_3_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_3_BYTE_OFFSET = 13'h0730;
  localparam int LDPC_DEC_EXPSYND_3_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_3_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_3_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_3_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_3_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_3_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_3_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_3_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_3_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_4_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_4_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_4_BYTE_OFFSET = 13'h0734;
  localparam int LDPC_DEC_EXPSYND_4_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_4_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_4_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_4_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_4_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_4_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_4_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_4_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_4_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_5_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_5_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_5_BYTE_OFFSET = 13'h0738;
  localparam int LDPC_DEC_EXPSYND_5_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_5_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_5_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_5_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_5_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_5_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_5_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_5_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_5_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_6_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_6_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_6_BYTE_OFFSET = 13'h073c;
  localparam int LDPC_DEC_EXPSYND_6_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_6_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_6_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_6_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_6_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_6_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_6_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_6_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_6_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_7_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_7_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_7_BYTE_OFFSET = 13'h0740;
  localparam int LDPC_DEC_EXPSYND_7_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_7_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_7_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_7_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_7_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_7_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_7_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_7_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_7_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_8_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_8_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_8_BYTE_OFFSET = 13'h0744;
  localparam int LDPC_DEC_EXPSYND_8_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_8_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_8_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_8_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_8_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_8_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_8_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_8_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_8_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_9_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_9_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_9_BYTE_OFFSET = 13'h0748;
  localparam int LDPC_DEC_EXPSYND_9_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_9_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_9_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_9_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_9_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_9_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_9_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_9_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_9_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_10_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_10_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_10_BYTE_OFFSET = 13'h074c;
  localparam int LDPC_DEC_EXPSYND_10_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_10_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_10_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_10_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_10_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_10_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_10_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_10_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_10_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_11_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_11_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_11_BYTE_OFFSET = 13'h0750;
  localparam int LDPC_DEC_EXPSYND_11_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_11_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_11_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_11_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_11_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_11_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_11_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_11_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_11_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_12_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_12_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_12_BYTE_OFFSET = 13'h0754;
  localparam int LDPC_DEC_EXPSYND_12_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_12_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_12_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_12_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_12_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_12_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_12_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_12_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_12_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_13_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_13_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_13_BYTE_OFFSET = 13'h0758;
  localparam int LDPC_DEC_EXPSYND_13_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_13_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_13_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_13_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_13_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_13_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_13_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_13_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_13_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_14_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_14_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_14_BYTE_OFFSET = 13'h075c;
  localparam int LDPC_DEC_EXPSYND_14_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_14_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_14_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_14_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_14_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_14_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_14_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_14_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_14_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_15_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_15_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_15_BYTE_OFFSET = 13'h0760;
  localparam int LDPC_DEC_EXPSYND_15_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_15_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_15_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_15_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_15_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_15_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_15_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_15_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_15_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_16_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_16_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_16_BYTE_OFFSET = 13'h0764;
  localparam int LDPC_DEC_EXPSYND_16_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_16_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_16_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_16_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_16_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_16_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_16_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_16_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_16_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_17_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_17_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_17_BYTE_OFFSET = 13'h0768;
  localparam int LDPC_DEC_EXPSYND_17_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_17_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_17_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_17_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_17_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_17_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_17_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_17_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_17_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_18_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_18_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_18_BYTE_OFFSET = 13'h076c;
  localparam int LDPC_DEC_EXPSYND_18_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_18_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_18_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_18_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_18_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_18_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_18_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_18_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_18_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_19_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_19_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_19_BYTE_OFFSET = 13'h0770;
  localparam int LDPC_DEC_EXPSYND_19_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_19_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_19_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_19_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_19_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_19_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_19_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_19_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_19_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_20_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_20_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_20_BYTE_OFFSET = 13'h0774;
  localparam int LDPC_DEC_EXPSYND_20_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_20_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_20_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_20_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_20_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_20_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_20_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_20_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_20_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_21_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_21_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_21_BYTE_OFFSET = 13'h0778;
  localparam int LDPC_DEC_EXPSYND_21_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_21_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_21_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_21_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_21_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_21_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_21_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_21_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_21_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_22_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_22_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_22_BYTE_OFFSET = 13'h077c;
  localparam int LDPC_DEC_EXPSYND_22_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_22_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_22_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_22_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_22_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_22_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_22_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_22_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_22_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_23_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_23_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_23_BYTE_OFFSET = 13'h0780;
  localparam int LDPC_DEC_EXPSYND_23_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_23_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_23_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_23_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_23_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_23_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_23_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_23_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_23_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_24_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_24_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_24_BYTE_OFFSET = 13'h0784;
  localparam int LDPC_DEC_EXPSYND_24_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_24_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_24_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_24_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_24_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_24_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_24_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_24_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_24_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_25_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_25_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_25_BYTE_OFFSET = 13'h0788;
  localparam int LDPC_DEC_EXPSYND_25_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_25_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_25_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_25_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_25_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_25_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_25_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_25_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_25_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_26_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_26_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_26_BYTE_OFFSET = 13'h078c;
  localparam int LDPC_DEC_EXPSYND_26_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_26_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_26_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_26_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_26_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_26_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_26_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_26_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_26_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_27_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_27_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_27_BYTE_OFFSET = 13'h0790;
  localparam int LDPC_DEC_EXPSYND_27_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_27_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_27_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_27_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_27_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_27_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_27_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_27_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_27_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_28_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_28_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_28_BYTE_OFFSET = 13'h0794;
  localparam int LDPC_DEC_EXPSYND_28_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_28_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_28_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_28_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_28_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_28_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_28_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_28_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_28_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_29_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_29_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_29_BYTE_OFFSET = 13'h0798;
  localparam int LDPC_DEC_EXPSYND_29_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_29_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_29_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_29_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_29_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_29_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_29_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_29_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_29_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_30_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_30_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_30_BYTE_OFFSET = 13'h079c;
  localparam int LDPC_DEC_EXPSYND_30_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_30_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_30_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_30_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_30_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_30_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_30_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_30_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_30_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_31_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_31_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_31_BYTE_OFFSET = 13'h07a0;
  localparam int LDPC_DEC_EXPSYND_31_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_31_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_31_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_31_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_31_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_31_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_31_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_31_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_31_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_32_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_32_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_32_BYTE_OFFSET = 13'h07a4;
  localparam int LDPC_DEC_EXPSYND_32_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_32_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_32_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_32_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_32_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_32_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_32_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_32_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_32_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_33_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_33_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_33_BYTE_OFFSET = 13'h07a8;
  localparam int LDPC_DEC_EXPSYND_33_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_33_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_33_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_33_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_33_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_33_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_33_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_33_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_33_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_34_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_34_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_34_BYTE_OFFSET = 13'h07ac;
  localparam int LDPC_DEC_EXPSYND_34_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_34_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_34_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_34_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_34_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_34_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_34_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_34_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_34_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_35_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_35_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_35_BYTE_OFFSET = 13'h07b0;
  localparam int LDPC_DEC_EXPSYND_35_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_35_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_35_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_35_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_35_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_35_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_35_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_35_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_35_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_36_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_36_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_36_BYTE_OFFSET = 13'h07b4;
  localparam int LDPC_DEC_EXPSYND_36_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_36_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_36_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_36_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_36_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_36_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_36_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_36_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_36_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_37_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_37_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_37_BYTE_OFFSET = 13'h07b8;
  localparam int LDPC_DEC_EXPSYND_37_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_37_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_37_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_37_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_37_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_37_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_37_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_37_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_37_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_38_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_38_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_38_BYTE_OFFSET = 13'h07bc;
  localparam int LDPC_DEC_EXPSYND_38_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_38_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_38_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_38_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_38_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_38_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_38_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_38_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_38_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_39_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_39_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_39_BYTE_OFFSET = 13'h07c0;
  localparam int LDPC_DEC_EXPSYND_39_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_39_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_39_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_39_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_39_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_39_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_39_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_39_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_39_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_40_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_40_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_40_BYTE_OFFSET = 13'h07c4;
  localparam int LDPC_DEC_EXPSYND_40_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_40_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_40_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_40_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_40_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_40_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_40_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_40_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_40_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_41_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_41_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_41_BYTE_OFFSET = 13'h07c8;
  localparam int LDPC_DEC_EXPSYND_41_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_41_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_41_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_41_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_41_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_41_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_41_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_41_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_41_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_42_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_42_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_42_BYTE_OFFSET = 13'h07cc;
  localparam int LDPC_DEC_EXPSYND_42_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_42_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_42_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_42_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_42_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_42_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_42_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_42_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_42_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_43_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_43_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_43_BYTE_OFFSET = 13'h07d0;
  localparam int LDPC_DEC_EXPSYND_43_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_43_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_43_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_43_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_43_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_43_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_43_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_43_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_43_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_44_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_44_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_44_BYTE_OFFSET = 13'h07d4;
  localparam int LDPC_DEC_EXPSYND_44_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_44_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_44_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_44_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_44_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_44_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_44_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_44_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_44_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_45_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_45_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_45_BYTE_OFFSET = 13'h07d8;
  localparam int LDPC_DEC_EXPSYND_45_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_45_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_45_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_45_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_45_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_45_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_45_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_45_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_45_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_46_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_46_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_46_BYTE_OFFSET = 13'h07dc;
  localparam int LDPC_DEC_EXPSYND_46_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_46_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_46_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_46_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_46_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_46_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_46_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_46_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_46_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_47_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_47_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_47_BYTE_OFFSET = 13'h07e0;
  localparam int LDPC_DEC_EXPSYND_47_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_47_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_47_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_47_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_47_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_47_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_47_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_47_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_47_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_48_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_48_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_48_BYTE_OFFSET = 13'h07e4;
  localparam int LDPC_DEC_EXPSYND_48_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_48_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_48_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_48_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_48_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_48_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_48_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_48_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_48_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_49_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_49_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_49_BYTE_OFFSET = 13'h07e8;
  localparam int LDPC_DEC_EXPSYND_49_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_49_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_49_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_49_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_49_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_49_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_49_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_49_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_49_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_50_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_50_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_50_BYTE_OFFSET = 13'h07ec;
  localparam int LDPC_DEC_EXPSYND_50_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_50_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_50_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_50_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_50_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_50_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_50_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_50_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_50_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_51_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_51_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_51_BYTE_OFFSET = 13'h07f0;
  localparam int LDPC_DEC_EXPSYND_51_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_51_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_51_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_51_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_51_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_51_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_51_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_51_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_51_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_52_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_52_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_52_BYTE_OFFSET = 13'h07f4;
  localparam int LDPC_DEC_EXPSYND_52_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_52_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_52_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_52_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_52_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_52_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_52_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_52_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_52_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_53_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_53_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_53_BYTE_OFFSET = 13'h07f8;
  localparam int LDPC_DEC_EXPSYND_53_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_53_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_53_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_53_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_53_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_53_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_53_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_53_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_53_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_54_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_54_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_54_BYTE_OFFSET = 13'h07fc;
  localparam int LDPC_DEC_EXPSYND_54_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_54_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_54_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_54_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_54_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_54_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_54_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_54_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_54_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_55_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_55_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_55_BYTE_OFFSET = 13'h0800;
  localparam int LDPC_DEC_EXPSYND_55_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_55_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_55_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_55_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_55_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_55_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_55_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_55_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_55_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_56_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_56_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_56_BYTE_OFFSET = 13'h0804;
  localparam int LDPC_DEC_EXPSYND_56_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_56_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_56_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_56_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_56_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_56_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_56_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_56_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_56_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_57_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_57_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_57_BYTE_OFFSET = 13'h0808;
  localparam int LDPC_DEC_EXPSYND_57_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_57_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_57_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_57_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_57_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_57_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_57_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_57_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_57_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_58_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_58_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_58_BYTE_OFFSET = 13'h080c;
  localparam int LDPC_DEC_EXPSYND_58_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_58_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_58_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_58_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_58_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_58_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_58_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_58_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_58_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_59_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_59_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_59_BYTE_OFFSET = 13'h0810;
  localparam int LDPC_DEC_EXPSYND_59_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_59_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_59_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_59_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_59_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_59_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_59_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_59_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_59_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_60_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_60_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_60_BYTE_OFFSET = 13'h0814;
  localparam int LDPC_DEC_EXPSYND_60_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_60_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_60_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_60_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_60_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_60_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_60_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_60_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_60_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_61_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_61_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_61_BYTE_OFFSET = 13'h0818;
  localparam int LDPC_DEC_EXPSYND_61_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_61_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_61_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_61_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_61_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_61_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_61_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_61_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_61_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_62_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_62_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_62_BYTE_OFFSET = 13'h081c;
  localparam int LDPC_DEC_EXPSYND_62_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_62_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_62_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_62_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_62_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_62_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_62_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_62_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_62_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_63_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_63_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_63_BYTE_OFFSET = 13'h0820;
  localparam int LDPC_DEC_EXPSYND_63_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_63_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_63_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_63_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_63_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_63_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_63_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_63_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_63_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_64_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_64_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_64_BYTE_OFFSET = 13'h0824;
  localparam int LDPC_DEC_EXPSYND_64_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_64_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_64_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_64_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_64_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_64_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_64_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_64_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_64_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_65_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_65_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_65_BYTE_OFFSET = 13'h0828;
  localparam int LDPC_DEC_EXPSYND_65_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_65_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_65_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_65_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_65_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_65_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_65_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_65_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_65_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_66_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_66_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_66_BYTE_OFFSET = 13'h082c;
  localparam int LDPC_DEC_EXPSYND_66_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_66_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_66_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_66_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_66_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_66_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_66_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_66_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_66_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_67_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_67_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_67_BYTE_OFFSET = 13'h0830;
  localparam int LDPC_DEC_EXPSYND_67_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_67_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_67_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_67_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_67_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_67_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_67_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_67_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_67_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_68_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_68_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_68_BYTE_OFFSET = 13'h0834;
  localparam int LDPC_DEC_EXPSYND_68_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_68_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_68_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_68_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_68_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_68_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_68_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_68_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_68_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_69_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_69_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_69_BYTE_OFFSET = 13'h0838;
  localparam int LDPC_DEC_EXPSYND_69_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_69_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_69_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_69_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_69_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_69_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_69_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_69_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_69_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_70_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_70_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_70_BYTE_OFFSET = 13'h083c;
  localparam int LDPC_DEC_EXPSYND_70_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_70_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_70_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_70_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_70_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_70_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_70_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_70_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_70_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_71_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_71_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_71_BYTE_OFFSET = 13'h0840;
  localparam int LDPC_DEC_EXPSYND_71_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_71_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_71_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_71_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_71_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_71_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_71_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_71_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_71_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_72_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_72_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_72_BYTE_OFFSET = 13'h0844;
  localparam int LDPC_DEC_EXPSYND_72_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_72_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_72_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_72_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_72_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_72_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_72_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_72_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_72_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_73_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_73_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_73_BYTE_OFFSET = 13'h0848;
  localparam int LDPC_DEC_EXPSYND_73_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_73_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_73_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_73_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_73_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_73_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_73_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_73_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_73_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_74_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_74_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_74_BYTE_OFFSET = 13'h084c;
  localparam int LDPC_DEC_EXPSYND_74_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_74_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_74_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_74_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_74_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_74_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_74_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_74_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_74_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_75_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_75_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_75_BYTE_OFFSET = 13'h0850;
  localparam int LDPC_DEC_EXPSYND_75_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_75_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_75_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_75_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_75_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_75_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_75_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_75_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_75_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_76_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_76_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_76_BYTE_OFFSET = 13'h0854;
  localparam int LDPC_DEC_EXPSYND_76_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_76_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_76_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_76_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_76_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_76_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_76_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_76_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_76_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_77_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_77_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_77_BYTE_OFFSET = 13'h0858;
  localparam int LDPC_DEC_EXPSYND_77_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_77_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_77_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_77_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_77_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_77_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_77_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_77_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_77_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_78_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_78_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_78_BYTE_OFFSET = 13'h085c;
  localparam int LDPC_DEC_EXPSYND_78_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_78_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_78_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_78_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_78_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_78_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_78_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_78_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_78_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_79_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_79_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_79_BYTE_OFFSET = 13'h0860;
  localparam int LDPC_DEC_EXPSYND_79_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_79_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_79_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_79_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_79_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_79_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_79_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_79_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_79_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_80_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_80_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_80_BYTE_OFFSET = 13'h0864;
  localparam int LDPC_DEC_EXPSYND_80_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_80_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_80_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_80_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_80_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_80_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_80_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_80_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_80_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_81_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_81_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_81_BYTE_OFFSET = 13'h0868;
  localparam int LDPC_DEC_EXPSYND_81_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_81_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_81_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_81_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_81_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_81_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_81_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_81_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_81_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_82_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_82_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_82_BYTE_OFFSET = 13'h086c;
  localparam int LDPC_DEC_EXPSYND_82_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_82_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_82_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_82_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_82_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_82_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_82_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_82_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_82_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_83_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_83_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_83_BYTE_OFFSET = 13'h0870;
  localparam int LDPC_DEC_EXPSYND_83_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_83_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_83_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_83_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_83_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_83_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_83_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_83_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_83_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_84_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_84_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_84_BYTE_OFFSET = 13'h0874;
  localparam int LDPC_DEC_EXPSYND_84_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_84_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_84_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_84_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_84_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_84_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_84_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_84_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_84_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_85_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_85_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_85_BYTE_OFFSET = 13'h0878;
  localparam int LDPC_DEC_EXPSYND_85_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_85_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_85_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_85_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_85_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_85_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_85_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_85_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_85_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_86_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_86_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_86_BYTE_OFFSET = 13'h087c;
  localparam int LDPC_DEC_EXPSYND_86_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_86_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_86_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_86_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_86_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_86_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_86_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_86_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_86_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_87_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_87_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_87_BYTE_OFFSET = 13'h0880;
  localparam int LDPC_DEC_EXPSYND_87_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_87_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_87_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_87_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_87_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_87_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_87_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_87_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_87_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_88_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_88_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_88_BYTE_OFFSET = 13'h0884;
  localparam int LDPC_DEC_EXPSYND_88_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_88_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_88_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_88_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_88_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_88_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_88_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_88_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_88_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_89_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_89_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_89_BYTE_OFFSET = 13'h0888;
  localparam int LDPC_DEC_EXPSYND_89_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_89_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_89_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_89_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_89_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_89_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_89_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_89_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_89_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_90_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_90_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_90_BYTE_OFFSET = 13'h088c;
  localparam int LDPC_DEC_EXPSYND_90_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_90_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_90_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_90_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_90_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_90_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_90_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_90_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_90_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_91_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_91_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_91_BYTE_OFFSET = 13'h0890;
  localparam int LDPC_DEC_EXPSYND_91_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_91_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_91_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_91_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_91_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_91_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_91_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_91_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_91_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_92_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_92_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_92_BYTE_OFFSET = 13'h0894;
  localparam int LDPC_DEC_EXPSYND_92_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_92_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_92_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_92_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_92_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_92_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_92_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_92_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_92_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_93_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_93_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_93_BYTE_OFFSET = 13'h0898;
  localparam int LDPC_DEC_EXPSYND_93_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_93_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_93_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_93_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_93_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_93_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_93_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_93_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_93_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_94_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_94_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_94_BYTE_OFFSET = 13'h089c;
  localparam int LDPC_DEC_EXPSYND_94_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_94_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_94_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_94_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_94_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_94_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_94_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_94_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_94_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_95_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_95_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_95_BYTE_OFFSET = 13'h08a0;
  localparam int LDPC_DEC_EXPSYND_95_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_95_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_95_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_95_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_95_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_95_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_95_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_95_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_95_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_96_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_96_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_96_BYTE_OFFSET = 13'h08a4;
  localparam int LDPC_DEC_EXPSYND_96_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_96_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_96_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_96_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_96_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_96_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_96_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_96_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_96_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_97_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_97_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_97_BYTE_OFFSET = 13'h08a8;
  localparam int LDPC_DEC_EXPSYND_97_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_97_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_97_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_97_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_97_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_97_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_97_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_97_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_97_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_98_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_98_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_98_BYTE_OFFSET = 13'h08ac;
  localparam int LDPC_DEC_EXPSYND_98_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_98_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_98_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_98_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_98_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_98_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_98_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_98_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_98_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_99_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_99_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_99_BYTE_OFFSET = 13'h08b0;
  localparam int LDPC_DEC_EXPSYND_99_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_99_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_99_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_99_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_99_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_99_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_99_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_99_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_99_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_100_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_100_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_100_BYTE_OFFSET = 13'h08b4;
  localparam int LDPC_DEC_EXPSYND_100_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_100_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_100_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_100_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_100_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_100_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_100_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_100_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_100_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_101_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_101_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_101_BYTE_OFFSET = 13'h08b8;
  localparam int LDPC_DEC_EXPSYND_101_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_101_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_101_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_101_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_101_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_101_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_101_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_101_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_101_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_102_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_102_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_102_BYTE_OFFSET = 13'h08bc;
  localparam int LDPC_DEC_EXPSYND_102_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_102_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_102_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_102_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_102_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_102_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_102_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_102_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_102_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_103_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_103_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_103_BYTE_OFFSET = 13'h08c0;
  localparam int LDPC_DEC_EXPSYND_103_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_103_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_103_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_103_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_103_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_103_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_103_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_103_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_103_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_104_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_104_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_104_BYTE_OFFSET = 13'h08c4;
  localparam int LDPC_DEC_EXPSYND_104_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_104_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_104_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_104_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_104_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_104_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_104_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_104_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_104_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_105_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_105_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_105_BYTE_OFFSET = 13'h08c8;
  localparam int LDPC_DEC_EXPSYND_105_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_105_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_105_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_105_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_105_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_105_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_105_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_105_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_105_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_106_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_106_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_106_BYTE_OFFSET = 13'h08cc;
  localparam int LDPC_DEC_EXPSYND_106_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_106_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_106_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_106_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_106_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_106_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_106_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_106_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_106_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_107_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_107_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_107_BYTE_OFFSET = 13'h08d0;
  localparam int LDPC_DEC_EXPSYND_107_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_107_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_107_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_107_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_107_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_107_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_107_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_107_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_107_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_108_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_108_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_108_BYTE_OFFSET = 13'h08d4;
  localparam int LDPC_DEC_EXPSYND_108_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_108_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_108_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_108_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_108_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_108_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_108_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_108_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_108_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_109_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_109_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_109_BYTE_OFFSET = 13'h08d8;
  localparam int LDPC_DEC_EXPSYND_109_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_109_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_109_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_109_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_109_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_109_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_109_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_109_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_109_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_110_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_110_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_110_BYTE_OFFSET = 13'h08dc;
  localparam int LDPC_DEC_EXPSYND_110_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_110_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_110_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_110_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_110_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_110_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_110_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_110_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_110_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_111_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_111_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_111_BYTE_OFFSET = 13'h08e0;
  localparam int LDPC_DEC_EXPSYND_111_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_111_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_111_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_111_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_111_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_111_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_111_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_111_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_111_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_112_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_112_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_112_BYTE_OFFSET = 13'h08e4;
  localparam int LDPC_DEC_EXPSYND_112_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_112_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_112_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_112_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_112_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_112_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_112_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_112_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_112_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_113_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_113_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_113_BYTE_OFFSET = 13'h08e8;
  localparam int LDPC_DEC_EXPSYND_113_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_113_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_113_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_113_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_113_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_113_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_113_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_113_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_113_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_114_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_114_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_114_BYTE_OFFSET = 13'h08ec;
  localparam int LDPC_DEC_EXPSYND_114_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_114_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_114_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_114_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_114_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_114_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_114_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_114_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_114_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_115_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_115_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_115_BYTE_OFFSET = 13'h08f0;
  localparam int LDPC_DEC_EXPSYND_115_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_115_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_115_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_115_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_115_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_115_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_115_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_115_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_115_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_116_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_116_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_116_BYTE_OFFSET = 13'h08f4;
  localparam int LDPC_DEC_EXPSYND_116_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_116_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_116_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_116_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_116_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_116_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_116_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_116_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_116_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_117_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_117_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_117_BYTE_OFFSET = 13'h08f8;
  localparam int LDPC_DEC_EXPSYND_117_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_117_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_117_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_117_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_117_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_117_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_117_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_117_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_117_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_118_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_118_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_118_BYTE_OFFSET = 13'h08fc;
  localparam int LDPC_DEC_EXPSYND_118_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_118_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_118_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_118_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_118_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_118_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_118_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_118_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_118_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_119_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_119_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_119_BYTE_OFFSET = 13'h0900;
  localparam int LDPC_DEC_EXPSYND_119_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_119_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_119_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_119_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_119_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_119_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_119_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_119_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_119_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_120_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_120_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_120_BYTE_OFFSET = 13'h0904;
  localparam int LDPC_DEC_EXPSYND_120_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_120_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_120_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_120_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_120_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_120_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_120_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_120_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_120_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_121_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_121_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_121_BYTE_OFFSET = 13'h0908;
  localparam int LDPC_DEC_EXPSYND_121_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_121_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_121_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_121_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_121_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_121_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_121_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_121_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_121_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_122_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_122_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_122_BYTE_OFFSET = 13'h090c;
  localparam int LDPC_DEC_EXPSYND_122_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_122_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_122_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_122_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_122_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_122_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_122_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_122_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_122_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_123_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_123_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_123_BYTE_OFFSET = 13'h0910;
  localparam int LDPC_DEC_EXPSYND_123_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_123_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_123_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_123_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_123_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_123_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_123_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_123_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_123_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_124_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_124_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_124_BYTE_OFFSET = 13'h0914;
  localparam int LDPC_DEC_EXPSYND_124_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_124_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_124_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_124_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_124_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_124_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_124_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_124_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_124_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_125_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_125_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_125_BYTE_OFFSET = 13'h0918;
  localparam int LDPC_DEC_EXPSYND_125_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_125_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_125_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_125_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_125_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_125_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_125_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_125_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_125_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_126_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_126_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_126_BYTE_OFFSET = 13'h091c;
  localparam int LDPC_DEC_EXPSYND_126_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_126_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_126_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_126_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_126_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_126_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_126_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_126_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_126_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_127_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_127_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_127_BYTE_OFFSET = 13'h0920;
  localparam int LDPC_DEC_EXPSYND_127_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_127_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_127_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_127_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_127_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_127_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_127_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_127_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_127_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_128_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_128_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_128_BYTE_OFFSET = 13'h0924;
  localparam int LDPC_DEC_EXPSYND_128_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_128_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_128_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_128_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_128_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_128_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_128_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_128_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_128_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_129_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_129_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_129_BYTE_OFFSET = 13'h0928;
  localparam int LDPC_DEC_EXPSYND_129_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_129_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_129_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_129_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_129_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_129_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_129_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_129_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_129_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_130_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_130_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_130_BYTE_OFFSET = 13'h092c;
  localparam int LDPC_DEC_EXPSYND_130_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_130_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_130_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_130_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_130_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_130_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_130_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_130_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_130_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_131_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_131_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_131_BYTE_OFFSET = 13'h0930;
  localparam int LDPC_DEC_EXPSYND_131_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_131_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_131_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_131_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_131_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_131_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_131_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_131_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_131_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_132_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_132_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_132_BYTE_OFFSET = 13'h0934;
  localparam int LDPC_DEC_EXPSYND_132_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_132_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_132_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_132_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_132_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_132_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_132_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_132_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_132_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_133_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_133_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_133_BYTE_OFFSET = 13'h0938;
  localparam int LDPC_DEC_EXPSYND_133_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_133_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_133_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_133_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_133_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_133_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_133_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_133_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_133_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_134_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_134_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_134_BYTE_OFFSET = 13'h093c;
  localparam int LDPC_DEC_EXPSYND_134_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_134_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_134_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_134_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_134_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_134_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_134_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_134_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_134_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_135_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_135_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_135_BYTE_OFFSET = 13'h0940;
  localparam int LDPC_DEC_EXPSYND_135_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_135_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_135_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_135_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_135_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_135_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_135_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_135_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_135_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_136_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_136_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_136_BYTE_OFFSET = 13'h0944;
  localparam int LDPC_DEC_EXPSYND_136_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_136_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_136_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_136_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_136_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_136_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_136_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_136_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_136_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_137_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_137_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_137_BYTE_OFFSET = 13'h0948;
  localparam int LDPC_DEC_EXPSYND_137_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_137_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_137_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_137_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_137_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_137_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_137_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_137_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_137_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_138_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_138_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_138_BYTE_OFFSET = 13'h094c;
  localparam int LDPC_DEC_EXPSYND_138_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_138_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_138_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_138_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_138_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_138_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_138_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_138_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_138_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_139_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_139_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_139_BYTE_OFFSET = 13'h0950;
  localparam int LDPC_DEC_EXPSYND_139_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_139_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_139_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_139_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_139_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_139_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_139_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_139_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_139_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_140_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_140_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_140_BYTE_OFFSET = 13'h0954;
  localparam int LDPC_DEC_EXPSYND_140_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_140_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_140_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_140_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_140_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_140_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_140_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_140_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_140_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_141_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_141_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_141_BYTE_OFFSET = 13'h0958;
  localparam int LDPC_DEC_EXPSYND_141_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_141_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_141_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_141_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_141_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_141_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_141_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_141_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_141_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_142_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_142_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_142_BYTE_OFFSET = 13'h095c;
  localparam int LDPC_DEC_EXPSYND_142_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_142_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_142_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_142_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_142_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_142_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_142_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_142_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_142_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_143_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_143_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_143_BYTE_OFFSET = 13'h0960;
  localparam int LDPC_DEC_EXPSYND_143_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_143_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_143_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_143_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_143_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_143_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_143_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_143_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_143_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_144_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_144_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_144_BYTE_OFFSET = 13'h0964;
  localparam int LDPC_DEC_EXPSYND_144_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_144_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_144_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_144_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_144_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_144_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_144_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_144_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_144_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_145_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_145_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_145_BYTE_OFFSET = 13'h0968;
  localparam int LDPC_DEC_EXPSYND_145_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_145_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_145_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_145_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_145_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_145_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_145_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_145_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_145_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_146_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_146_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_146_BYTE_OFFSET = 13'h096c;
  localparam int LDPC_DEC_EXPSYND_146_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_146_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_146_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_146_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_146_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_146_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_146_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_146_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_146_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_147_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_147_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_147_BYTE_OFFSET = 13'h0970;
  localparam int LDPC_DEC_EXPSYND_147_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_147_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_147_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_147_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_147_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_147_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_147_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_147_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_147_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_148_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_148_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_148_BYTE_OFFSET = 13'h0974;
  localparam int LDPC_DEC_EXPSYND_148_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_148_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_148_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_148_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_148_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_148_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_148_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_148_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_148_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_149_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_149_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_149_BYTE_OFFSET = 13'h0978;
  localparam int LDPC_DEC_EXPSYND_149_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_149_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_149_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_149_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_149_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_149_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_149_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_149_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_149_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_150_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_150_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_150_BYTE_OFFSET = 13'h097c;
  localparam int LDPC_DEC_EXPSYND_150_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_150_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_150_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_150_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_150_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_150_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_150_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_150_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_150_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_151_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_151_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_151_BYTE_OFFSET = 13'h0980;
  localparam int LDPC_DEC_EXPSYND_151_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_151_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_151_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_151_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_151_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_151_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_151_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_151_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_151_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_152_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_152_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_152_BYTE_OFFSET = 13'h0984;
  localparam int LDPC_DEC_EXPSYND_152_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_152_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_152_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_152_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_152_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_152_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_152_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_152_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_152_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_153_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_153_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_153_BYTE_OFFSET = 13'h0988;
  localparam int LDPC_DEC_EXPSYND_153_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_153_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_153_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_153_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_153_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_153_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_153_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_153_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_153_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_154_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_154_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_154_BYTE_OFFSET = 13'h098c;
  localparam int LDPC_DEC_EXPSYND_154_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_154_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_154_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_154_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_154_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_154_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_154_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_154_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_154_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_155_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_155_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_155_BYTE_OFFSET = 13'h0990;
  localparam int LDPC_DEC_EXPSYND_155_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_155_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_155_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_155_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_155_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_155_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_155_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_155_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_155_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_156_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_156_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_156_BYTE_OFFSET = 13'h0994;
  localparam int LDPC_DEC_EXPSYND_156_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_156_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_156_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_156_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_156_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_156_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_156_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_156_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_156_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_157_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_157_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_157_BYTE_OFFSET = 13'h0998;
  localparam int LDPC_DEC_EXPSYND_157_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_157_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_157_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_157_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_157_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_157_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_157_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_157_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_157_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_158_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_158_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_158_BYTE_OFFSET = 13'h099c;
  localparam int LDPC_DEC_EXPSYND_158_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_158_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_158_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_158_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_158_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_158_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_158_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_158_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_158_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_159_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_159_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_159_BYTE_OFFSET = 13'h09a0;
  localparam int LDPC_DEC_EXPSYND_159_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_159_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_159_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_159_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_159_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_159_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_159_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_159_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_159_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_160_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_160_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_160_BYTE_OFFSET = 13'h09a4;
  localparam int LDPC_DEC_EXPSYND_160_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_160_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_160_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_160_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_160_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_160_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_160_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_160_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_160_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_161_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_161_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_161_BYTE_OFFSET = 13'h09a8;
  localparam int LDPC_DEC_EXPSYND_161_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_161_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_161_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_161_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_161_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_161_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_161_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_161_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_161_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_162_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_162_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_162_BYTE_OFFSET = 13'h09ac;
  localparam int LDPC_DEC_EXPSYND_162_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_162_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_162_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_162_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_162_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_162_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_162_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_162_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_162_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_163_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_163_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_163_BYTE_OFFSET = 13'h09b0;
  localparam int LDPC_DEC_EXPSYND_163_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_163_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_163_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_163_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_163_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_163_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_163_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_163_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_163_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_164_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_164_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_164_BYTE_OFFSET = 13'h09b4;
  localparam int LDPC_DEC_EXPSYND_164_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_164_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_164_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_164_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_164_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_164_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_164_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_164_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_164_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_165_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_165_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_165_BYTE_OFFSET = 13'h09b8;
  localparam int LDPC_DEC_EXPSYND_165_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_165_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_165_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_165_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_165_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_165_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_165_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_165_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_165_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_166_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_166_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_166_BYTE_OFFSET = 13'h09bc;
  localparam int LDPC_DEC_EXPSYND_166_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_166_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_166_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_166_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_166_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_166_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_166_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_166_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_166_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_EXPSYND_167_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_167_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_167_BYTE_OFFSET = 13'h09c0;
  localparam int LDPC_DEC_EXPSYND_167_EXP_SYNR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_167_EXP_SYNR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_167_EXP_SYNR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_167_EXP_SYNW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_167_EXP_SYNW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_167_EXP_SYNW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_EXPSYND_167_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_EXPSYND_167_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_EXPSYND_167_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_PROBABILITY_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_PROBABILITY_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_PROBABILITY_BYTE_OFFSET = 13'h09c4;
  localparam int LDPC_DEC_PROBABILITY_PERC_PROBABILITY_BIT_WIDTH = 32;
  localparam bit [31:0] LDPC_DEC_PROBABILITY_PERC_PROBABILITY_BIT_MASK = 32'hffffffff;
  localparam int LDPC_DEC_PROBABILITY_PERC_PROBABILITY_BIT_OFFSET = 0;
  localparam int LDPC_DEC_HAMDIST_LOOP_MAX_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_HAMDIST_LOOP_MAX_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_HAMDIST_LOOP_MAX_BYTE_OFFSET = 13'h09c8;
  localparam int LDPC_DEC_HAMDIST_LOOP_MAX_HAMDIST_LOOP_MAX_BIT_WIDTH = 32;
  localparam bit [31:0] LDPC_DEC_HAMDIST_LOOP_MAX_HAMDIST_LOOP_MAX_BIT_MASK = 32'hffffffff;
  localparam int LDPC_DEC_HAMDIST_LOOP_MAX_HAMDIST_LOOP_MAX_BIT_OFFSET = 0;
  localparam int LDPC_DEC_HAMDIST_LOOP_PERCENTAGE_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_HAMDIST_LOOP_PERCENTAGE_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_HAMDIST_LOOP_PERCENTAGE_BYTE_OFFSET = 13'h09cc;
  localparam int LDPC_DEC_HAMDIST_LOOP_PERCENTAGE_HAMDIST_LOOP_PERCENTAGE_BIT_WIDTH = 32;
  localparam bit [31:0] LDPC_DEC_HAMDIST_LOOP_PERCENTAGE_HAMDIST_LOOP_PERCENTAGE_BIT_MASK = 32'hffffffff;
  localparam int LDPC_DEC_HAMDIST_LOOP_PERCENTAGE_HAMDIST_LOOP_PERCENTAGE_BIT_OFFSET = 0;
  localparam int LDPC_DEC_HAMDIST_IIR1_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_HAMDIST_IIR1_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_HAMDIST_IIR1_BYTE_OFFSET = 13'h09d0;
  localparam int LDPC_DEC_HAMDIST_IIR1_HAMDIST_IIR1_BIT_WIDTH = 32;
  localparam bit [31:0] LDPC_DEC_HAMDIST_IIR1_HAMDIST_IIR1_BIT_MASK = 32'hffffffff;
  localparam int LDPC_DEC_HAMDIST_IIR1_HAMDIST_IIR1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_HAMDIST_IIR2_NOT_USED_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_HAMDIST_IIR2_NOT_USED_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_HAMDIST_IIR2_NOT_USED_BYTE_OFFSET = 13'h09d4;
  localparam int LDPC_DEC_HAMDIST_IIR2_NOT_USED_HAMDIST_IIR2_BIT_WIDTH = 32;
  localparam bit [31:0] LDPC_DEC_HAMDIST_IIR2_NOT_USED_HAMDIST_IIR2_BIT_MASK = 32'hffffffff;
  localparam int LDPC_DEC_HAMDIST_IIR2_NOT_USED_HAMDIST_IIR2_BIT_OFFSET = 0;
  localparam int LDPC_DEC_HAMDIST_IIR3_NOT_USED_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_HAMDIST_IIR3_NOT_USED_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_HAMDIST_IIR3_NOT_USED_BYTE_OFFSET = 13'h09d8;
  localparam int LDPC_DEC_HAMDIST_IIR3_NOT_USED_HAMDIST_IIR3_BIT_WIDTH = 32;
  localparam bit [31:0] LDPC_DEC_HAMDIST_IIR3_NOT_USED_HAMDIST_IIR3_BIT_MASK = 32'hffffffff;
  localparam int LDPC_DEC_HAMDIST_IIR3_NOT_USED_HAMDIST_IIR3_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CONVERGED_VALID_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CONVERGED_VALID_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CONVERGED_VALID_BYTE_OFFSET = 13'h09dc;
  localparam int LDPC_DEC_CONVERGED_VALID_CONVERGEDR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CONVERGED_VALID_CONVERGEDR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CONVERGED_VALID_CONVERGEDR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CONVERGED_VALID_CONVERGEDW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CONVERGED_VALID_CONVERGEDW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CONVERGED_VALID_CONVERGEDW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_CONVERGED_VALID_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_CONVERGED_VALID_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_CONVERGED_VALID_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CONVERGED_STATUS_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CONVERGED_STATUS_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CONVERGED_STATUS_BYTE_OFFSET = 13'h09e0;
  localparam int LDPC_DEC_CONVERGED_STATUS_CONVERGEDR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CONVERGED_STATUS_CONVERGEDR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CONVERGED_STATUS_CONVERGEDR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CONVERGED_STATUS_CONVERGEDW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CONVERGED_STATUS_CONVERGEDW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CONVERGED_STATUS_CONVERGEDW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_CONVERGED_STATUS_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_CONVERGED_STATUS_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_CONVERGED_STATUS_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_CONVERGED_VALID_NOT_USED_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CONVERGED_VALID_NOT_USED_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CONVERGED_VALID_NOT_USED_BYTE_OFFSET = 13'h09e4;
  localparam int LDPC_DEC_CONVERGED_VALID_NOT_USED_CONVERGED_VALIDR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CONVERGED_VALID_NOT_USED_CONVERGED_VALIDR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CONVERGED_VALID_NOT_USED_CONVERGED_VALIDR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CONVERGED_VALID_NOT_USED_CONVERGED_VALIDW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CONVERGED_VALID_NOT_USED_CONVERGED_VALIDW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CONVERGED_VALID_NOT_USED_CONVERGED_VALIDW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_CONVERGED_VALID_NOT_USED_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_CONVERGED_VALID_NOT_USED_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_CONVERGED_VALID_NOT_USED_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_START_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_START_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_START_BYTE_OFFSET = 13'h09e8;
  localparam int LDPC_DEC_START_STARTR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_START_STARTR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_START_STARTR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_START_STARTW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_START_STARTW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_START_STARTW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_START_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_START_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_START_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_VALID_NOT_USED_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_VALID_NOT_USED_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_VALID_NOT_USED_BYTE_OFFSET = 13'h09ec;
  localparam int LDPC_DEC_VALID_NOT_USED_VALIDR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_VALID_NOT_USED_VALIDR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_VALID_NOT_USED_VALIDR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_VALID_NOT_USED_VALIDW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_VALID_NOT_USED_VALIDW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_VALID_NOT_USED_VALIDW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_VALID_NOT_USED_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_VALID_NOT_USED_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_VALID_NOT_USED_RESERVED_BIT_OFFSET = 2;
  localparam int LDPC_DEC_VALID_CODEWORD_NOT_USED_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_VALID_CODEWORD_NOT_USED_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_VALID_CODEWORD_NOT_USED_BYTE_OFFSET = 13'h09f0;
  localparam int LDPC_DEC_VALID_CODEWORD_NOT_USED_VALID_CODEWORDR_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_VALID_CODEWORD_NOT_USED_VALID_CODEWORDR_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_VALID_CODEWORD_NOT_USED_VALID_CODEWORDR_BIT_OFFSET = 0;
  localparam int LDPC_DEC_VALID_CODEWORD_NOT_USED_VALID_CODEWORDW_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_VALID_CODEWORD_NOT_USED_VALID_CODEWORDW_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_VALID_CODEWORD_NOT_USED_VALID_CODEWORDW_BIT_OFFSET = 1;
  localparam int LDPC_DEC_VALID_CODEWORD_NOT_USED_RESERVED_BIT_WIDTH = 30;
  localparam bit [29:0] LDPC_DEC_VALID_CODEWORD_NOT_USED_RESERVED_BIT_MASK = 30'h3fffffff;
  localparam int LDPC_DEC_VALID_CODEWORD_NOT_USED_RESERVED_BIT_OFFSET = 2;
endpackage
