`include "GF2_LDPC_flogtanh_0x00000_inc.sv"
`include "GF2_LDPC_flogtanh_0x00001_inc.sv"
`include "GF2_LDPC_flogtanh_0x00002_inc.sv"
`include "GF2_LDPC_flogtanh_0x00003_inc.sv"
`include "GF2_LDPC_flogtanh_0x00004_inc.sv"
`include "GF2_LDPC_flogtanh_0x00005_inc.sv"
`include "GF2_LDPC_flogtanh_0x00006_inc.sv"
`include "GF2_LDPC_flogtanh_0x00007_inc.sv"
`include "GF2_LDPC_flogtanh_0x00008_inc.sv"
`include "GF2_LDPC_flogtanh_0x00009_inc.sv"
