              flogtanh0x00008_0 = 
          (!flogtanh_sel[7]) ? 
                       flogtanh0x00007_0_q: 
                       flogtanh0x00007_1_q;
              flogtanh0x00008_1 = 
          (!flogtanh_sel[7]) ? 
                       flogtanh0x00007_2_q: 
                       flogtanh0x00007_3_q;
