parameter MAX_SUM_WDTH = 11 ,
