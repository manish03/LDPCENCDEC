              fgallag0x00007_0 = 
          (!fgallag_sel[6]) ? 
                       fgallag0x00006_0_q: 
                       fgallag0x00006_1_q;
              fgallag0x00007_1 = 
          (!fgallag_sel[6]) ? 
                       fgallag0x00006_2_q: 
                       fgallag0x00006_3_q;
              fgallag0x00007_2 = 
          (!fgallag_sel[6]) ? 
                       fgallag0x00006_4_q: 
                       fgallag0x00006_5_q;
               fgallag0x00007_3 =  0;
