reg [flogtanh_WDTH -1:0] flogtanh0x00003_0, flogtanh0x00003_0_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00003_1, flogtanh0x00003_1_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00003_2, flogtanh0x00003_2_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00003_3, flogtanh0x00003_3_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00003_4, flogtanh0x00003_4_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00003_5, flogtanh0x00003_5_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00003_6, flogtanh0x00003_6_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00003_7, flogtanh0x00003_7_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00003_8, flogtanh0x00003_8_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00003_9, flogtanh0x00003_9_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00003_10, flogtanh0x00003_10_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00003_11, flogtanh0x00003_11_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00003_12, flogtanh0x00003_12_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00003_13, flogtanh0x00003_13_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00003_14, flogtanh0x00003_14_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00003_15, flogtanh0x00003_15_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00003_16, flogtanh0x00003_16_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00003_17, flogtanh0x00003_17_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00003_18, flogtanh0x00003_18_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00003_19, flogtanh0x00003_19_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00003_20, flogtanh0x00003_20_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00003_21, flogtanh0x00003_21_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00003_22, flogtanh0x00003_22_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00003_23, flogtanh0x00003_23_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00003_24, flogtanh0x00003_24_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00003_25, flogtanh0x00003_25_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00003_26, flogtanh0x00003_26_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00003_27, flogtanh0x00003_27_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00003_28, flogtanh0x00003_28_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00003_29, flogtanh0x00003_29_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00003_30, flogtanh0x00003_30_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00003_31, flogtanh0x00003_31_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00003_32, flogtanh0x00003_32_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00003_33, flogtanh0x00003_33_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00003_34, flogtanh0x00003_34_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00003_35, flogtanh0x00003_35_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00003_36, flogtanh0x00003_36_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00003_37, flogtanh0x00003_37_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00003_38, flogtanh0x00003_38_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00003_39, flogtanh0x00003_39_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00003_40, flogtanh0x00003_40_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00003_41, flogtanh0x00003_41_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00003_42, flogtanh0x00003_42_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00003_43, flogtanh0x00003_43_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00003_44, flogtanh0x00003_44_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00003_45, flogtanh0x00003_45_q;
reg start_d_flogtanh0x00003_q ;
always_comb begin
 flogtanh0x00003_0_q =  flogtanh0x00003_0;
 flogtanh0x00003_1_q =  flogtanh0x00003_1;
 flogtanh0x00003_2_q =  flogtanh0x00003_2;
 flogtanh0x00003_3_q =  flogtanh0x00003_3;
 flogtanh0x00003_4_q =  flogtanh0x00003_4;
 flogtanh0x00003_5_q =  flogtanh0x00003_5;
 flogtanh0x00003_6_q =  flogtanh0x00003_6;
 flogtanh0x00003_7_q =  flogtanh0x00003_7;
 flogtanh0x00003_8_q =  flogtanh0x00003_8;
 flogtanh0x00003_9_q =  flogtanh0x00003_9;
 flogtanh0x00003_10_q =  flogtanh0x00003_10;
 flogtanh0x00003_11_q =  flogtanh0x00003_11;
 flogtanh0x00003_12_q =  flogtanh0x00003_12;
 flogtanh0x00003_13_q =  flogtanh0x00003_13;
 flogtanh0x00003_14_q =  flogtanh0x00003_14;
 flogtanh0x00003_15_q =  flogtanh0x00003_15;
 flogtanh0x00003_16_q =  flogtanh0x00003_16;
 flogtanh0x00003_17_q =  flogtanh0x00003_17;
 flogtanh0x00003_18_q =  flogtanh0x00003_18;
 flogtanh0x00003_19_q =  flogtanh0x00003_19;
 flogtanh0x00003_20_q =  flogtanh0x00003_20;
 flogtanh0x00003_21_q =  flogtanh0x00003_21;
 flogtanh0x00003_22_q =  flogtanh0x00003_22;
 flogtanh0x00003_23_q =  flogtanh0x00003_23;
 flogtanh0x00003_24_q =  flogtanh0x00003_24;
 flogtanh0x00003_25_q =  flogtanh0x00003_25;
 flogtanh0x00003_26_q =  flogtanh0x00003_26;
 flogtanh0x00003_27_q =  flogtanh0x00003_27;
 flogtanh0x00003_28_q =  flogtanh0x00003_28;
 flogtanh0x00003_29_q =  flogtanh0x00003_29;
 flogtanh0x00003_30_q =  flogtanh0x00003_30;
 flogtanh0x00003_31_q =  flogtanh0x00003_31;
 flogtanh0x00003_32_q =  flogtanh0x00003_32;
 flogtanh0x00003_33_q =  flogtanh0x00003_33;
 flogtanh0x00003_34_q =  flogtanh0x00003_34;
 flogtanh0x00003_35_q =  flogtanh0x00003_35;
 flogtanh0x00003_36_q =  flogtanh0x00003_36;
 flogtanh0x00003_37_q =  flogtanh0x00003_37;
 flogtanh0x00003_38_q =  flogtanh0x00003_38;
 flogtanh0x00003_39_q =  flogtanh0x00003_39;
 flogtanh0x00003_40_q =  flogtanh0x00003_40;
 flogtanh0x00003_41_q =  flogtanh0x00003_41;
 flogtanh0x00003_42_q =  flogtanh0x00003_42;
 flogtanh0x00003_43_q =  flogtanh0x00003_43;
 flogtanh0x00003_44_q =  flogtanh0x00003_44;
 flogtanh0x00003_45_q =  flogtanh0x00003_45;
 start_d_flogtanh0x00003_q =  start_d_flogtanh0x00002_q;
end
