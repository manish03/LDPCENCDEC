              fgallag0x00008_0 = 
          (!fgallag_sel[7]) ? 
                       fgallag0x00007_0_q: 
                       fgallag0x00007_1_q;
              fgallag0x00008_1 = 
          (!fgallag_sel[7]) ? 
                       fgallag0x00007_2_q: 
                       fgallag0x00007_3_q;
