reg [flogtanh_WDTH -1:0] flogtanh0xffffffff_0, flogtanh0xffffffff_0_q;
reg [flogtanh_WDTH -1:0] flogtanh0xffffffff_1, flogtanh0xffffffff_1_q;
reg start_d_flogtanh0xffffffff_q ;
always_comb begin
 flogtanh0xffffffff_0_q =  flogtanh0xffffffff_0;
 flogtanh0xffffffff_1_q =  flogtanh0xffffffff_1;
 start_d_flogtanh0xffffffff_q =  start_d_flogtanh0x00008_q;
end
