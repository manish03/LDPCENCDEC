always_comb
begin
`include "GF2_LDPC_fgallag_0x00000.sv"
end
always_comb
begin
`include "GF2_LDPC_fgallag_0x00001.sv"
end
always_comb
begin
`include "GF2_LDPC_fgallag_0x00002.sv"
end
always_comb
begin
`include "GF2_LDPC_fgallag_0x00003.sv"
end
always_comb
begin
`include "GF2_LDPC_fgallag_0x00004.sv"
end
always_comb
begin
`include "GF2_LDPC_fgallag_0x00005.sv"
end
always_comb
begin
`include "GF2_LDPC_fgallag_0x00006.sv"
end
always_comb
begin
`include "GF2_LDPC_fgallag_0x00007.sv"
end
always_comb
begin
`include "GF2_LDPC_fgallag_0x00008.sv"
end
always_comb
begin
`include "GF2_LDPC_fgallag_0x00009.sv"
end
