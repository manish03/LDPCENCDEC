parameter n_minus_m = 'd40;
parameter n_int = 'd208;
parameter m_int = 'd168;



parameter z_int = 'd4;



wire y_nr_40_0;
assign y_nr_40_0 = 
        y_nr_enc[1] ^ 
        y_nr_enc[5] ^ 
        y_nr_enc[8] ^ 
0; ///1



wire y_nr_40_1;
assign y_nr_40_1 = 
        y_nr_enc[14] ^ 
        y_nr_enc[25] ^ 
        y_nr_enc[37] ^ 
0; ///1



wire y_nr_40_2;
assign y_nr_40_2 = 
        y_nr_enc[3] ^ 
        y_nr_enc[14] ^ 
        y_nr_enc[17] ^ 
0; ///1



wire y_nr_40_3;
assign y_nr_40_3 = 
        y_nr_enc[21] ^ 
        y_nr_enc[26] ^ 
        y_nr_enc[28] ^ 
0; ///1



wire y_nr_40_4;
assign y_nr_40_4 = 
        y_nr_enc[32] ^ 
        y_nr_enc[36] ^ 
        y_nr_enc[1] ^ 
0; ///1



wire y_nr_40_5;
assign y_nr_40_5 = 
        y_nr_enc[6] ^ 
        y_nr_enc[12] ^ 
        y_nr_enc[16] ^ 
0; ///1



wire y_nr_40_6;
assign y_nr_40_6 = 
        y_nr_enc[32] ^ 
        y_nr_enc[4] ^ 
        y_nr_enc[10] ^ 
0; ///1



wire y_nr_40_7;
assign y_nr_40_7 = 
        y_nr_enc[18] ^ 
        y_nr_enc[20] ^ 
        y_nr_enc[25] ^ 
0; ///1



wire y_nr_40_8;
assign y_nr_40_8 = 
        y_nr_enc[30] ^ 
        y_nr_enc[34] ^ 
        y_nr_enc[36] ^ 
0; ///1



    assign y_nr_p40 = 
y_nr_40_0 ^ 
y_nr_40_1 ^ 
y_nr_40_2 ^ 
y_nr_40_3 ^ 
y_nr_40_4 ^ 
y_nr_40_5 ^ 
y_nr_40_6 ^ 
y_nr_40_7 ^ 
y_nr_40_8 ^ 
0; ///3



wire y_nr_41_0;
assign y_nr_41_0 = 
        y_nr_enc[2] ^ 
        y_nr_enc[6] ^ 
        y_nr_enc[9] ^ 
0; ///1



wire y_nr_41_1;
assign y_nr_41_1 = 
        y_nr_enc[15] ^ 
        y_nr_enc[26] ^ 
        y_nr_enc[38] ^ 
0; ///1



wire y_nr_41_2;
assign y_nr_41_2 = 
        y_nr_enc[0] ^ 
        y_nr_enc[15] ^ 
        y_nr_enc[18] ^ 
0; ///1



wire y_nr_41_3;
assign y_nr_41_3 = 
        y_nr_enc[22] ^ 
        y_nr_enc[27] ^ 
        y_nr_enc[29] ^ 
0; ///1



wire y_nr_41_4;
assign y_nr_41_4 = 
        y_nr_enc[33] ^ 
        y_nr_enc[37] ^ 
        y_nr_enc[2] ^ 
0; ///1



wire y_nr_41_5;
assign y_nr_41_5 = 
        y_nr_enc[7] ^ 
        y_nr_enc[13] ^ 
        y_nr_enc[17] ^ 
0; ///1



wire y_nr_41_6;
assign y_nr_41_6 = 
        y_nr_enc[33] ^ 
        y_nr_enc[5] ^ 
        y_nr_enc[11] ^ 
0; ///1



wire y_nr_41_7;
assign y_nr_41_7 = 
        y_nr_enc[19] ^ 
        y_nr_enc[21] ^ 
        y_nr_enc[26] ^ 
0; ///1



wire y_nr_41_8;
assign y_nr_41_8 = 
        y_nr_enc[31] ^ 
        y_nr_enc[35] ^ 
        y_nr_enc[37] ^ 
0; ///1



    assign y_nr_p41 = 
y_nr_41_0 ^ 
y_nr_41_1 ^ 
y_nr_41_2 ^ 
y_nr_41_3 ^ 
y_nr_41_4 ^ 
y_nr_41_5 ^ 
y_nr_41_6 ^ 
y_nr_41_7 ^ 
y_nr_41_8 ^ 
0; ///3



wire y_nr_42_0;
assign y_nr_42_0 = 
        y_nr_enc[3] ^ 
        y_nr_enc[7] ^ 
        y_nr_enc[10] ^ 
0; ///1



wire y_nr_42_1;
assign y_nr_42_1 = 
        y_nr_enc[12] ^ 
        y_nr_enc[27] ^ 
        y_nr_enc[39] ^ 
0; ///1



wire y_nr_42_2;
assign y_nr_42_2 = 
        y_nr_enc[1] ^ 
        y_nr_enc[12] ^ 
        y_nr_enc[19] ^ 
0; ///1



wire y_nr_42_3;
assign y_nr_42_3 = 
        y_nr_enc[23] ^ 
        y_nr_enc[24] ^ 
        y_nr_enc[30] ^ 
0; ///1



wire y_nr_42_4;
assign y_nr_42_4 = 
        y_nr_enc[34] ^ 
        y_nr_enc[38] ^ 
        y_nr_enc[3] ^ 
0; ///1



wire y_nr_42_5;
assign y_nr_42_5 = 
        y_nr_enc[4] ^ 
        y_nr_enc[14] ^ 
        y_nr_enc[18] ^ 
0; ///1



wire y_nr_42_6;
assign y_nr_42_6 = 
        y_nr_enc[34] ^ 
        y_nr_enc[6] ^ 
        y_nr_enc[8] ^ 
0; ///1



wire y_nr_42_7;
assign y_nr_42_7 = 
        y_nr_enc[16] ^ 
        y_nr_enc[22] ^ 
        y_nr_enc[27] ^ 
0; ///1



wire y_nr_42_8;
assign y_nr_42_8 = 
        y_nr_enc[28] ^ 
        y_nr_enc[32] ^ 
        y_nr_enc[38] ^ 
0; ///1



    assign y_nr_p42 = 
y_nr_42_0 ^ 
y_nr_42_1 ^ 
y_nr_42_2 ^ 
y_nr_42_3 ^ 
y_nr_42_4 ^ 
y_nr_42_5 ^ 
y_nr_42_6 ^ 
y_nr_42_7 ^ 
y_nr_42_8 ^ 
0; ///3



wire y_nr_43_0;
assign y_nr_43_0 = 
        y_nr_enc[0] ^ 
        y_nr_enc[4] ^ 
        y_nr_enc[11] ^ 
0; ///1



wire y_nr_43_1;
assign y_nr_43_1 = 
        y_nr_enc[13] ^ 
        y_nr_enc[24] ^ 
        y_nr_enc[36] ^ 
0; ///1



wire y_nr_43_2;
assign y_nr_43_2 = 
        y_nr_enc[2] ^ 
        y_nr_enc[13] ^ 
        y_nr_enc[16] ^ 
0; ///1



wire y_nr_43_3;
assign y_nr_43_3 = 
        y_nr_enc[20] ^ 
        y_nr_enc[25] ^ 
        y_nr_enc[31] ^ 
0; ///1



wire y_nr_43_4;
assign y_nr_43_4 = 
        y_nr_enc[35] ^ 
        y_nr_enc[39] ^ 
        y_nr_enc[0] ^ 
0; ///1



wire y_nr_43_5;
assign y_nr_43_5 = 
        y_nr_enc[5] ^ 
        y_nr_enc[15] ^ 
        y_nr_enc[19] ^ 
0; ///1



wire y_nr_43_6;
assign y_nr_43_6 = 
        y_nr_enc[35] ^ 
        y_nr_enc[7] ^ 
        y_nr_enc[9] ^ 
0; ///1



wire y_nr_43_7;
assign y_nr_43_7 = 
        y_nr_enc[17] ^ 
        y_nr_enc[23] ^ 
        y_nr_enc[24] ^ 
0; ///1



wire y_nr_43_8;
assign y_nr_43_8 = 
        y_nr_enc[29] ^ 
        y_nr_enc[33] ^ 
        y_nr_enc[39] ^ 
0; ///1



    assign y_nr_p43 = 
y_nr_43_0 ^ 
y_nr_43_1 ^ 
y_nr_43_2 ^ 
y_nr_43_3 ^ 
y_nr_43_4 ^ 
y_nr_43_5 ^ 
y_nr_43_6 ^ 
y_nr_43_7 ^ 
y_nr_43_8 ^ 
0; ///3



wire y_nr_44_0;
assign y_nr_44_0 = 
        y_nr_enc[1] ^ 
        y_nr_enc[5] ^ 
        y_nr_enc[8] ^ 
0; ///1



wire y_nr_44_1;
assign y_nr_44_1 = 
        y_nr_enc[14] ^ 
        y_nr_enc[25] ^ 
        y_nr_enc[37] ^ 
0; ///1



wire y_nr_44_2;
assign y_nr_44_2 = 
        y_nr_enc[40] ^ 
0; ///1



    assign y_nr_p44 = 
y_nr_44_0 ^ 
y_nr_44_1 ^ 
y_nr_44_2 ^ 
0; ///3



wire y_nr_45_0;
assign y_nr_45_0 = 
        y_nr_enc[2] ^ 
        y_nr_enc[6] ^ 
        y_nr_enc[9] ^ 
0; ///1



wire y_nr_45_1;
assign y_nr_45_1 = 
        y_nr_enc[15] ^ 
        y_nr_enc[26] ^ 
        y_nr_enc[38] ^ 
0; ///1



wire y_nr_45_2;
assign y_nr_45_2 = 
        y_nr_enc[41] ^ 
0; ///1



    assign y_nr_p45 = 
y_nr_45_0 ^ 
y_nr_45_1 ^ 
y_nr_45_2 ^ 
0; ///3



wire y_nr_46_0;
assign y_nr_46_0 = 
        y_nr_enc[3] ^ 
        y_nr_enc[7] ^ 
        y_nr_enc[10] ^ 
0; ///1



wire y_nr_46_1;
assign y_nr_46_1 = 
        y_nr_enc[12] ^ 
        y_nr_enc[27] ^ 
        y_nr_enc[39] ^ 
0; ///1



wire y_nr_46_2;
assign y_nr_46_2 = 
        y_nr_enc[42] ^ 
0; ///1



    assign y_nr_p46 = 
y_nr_46_0 ^ 
y_nr_46_1 ^ 
y_nr_46_2 ^ 
0; ///3



wire y_nr_47_0;
assign y_nr_47_0 = 
        y_nr_enc[0] ^ 
        y_nr_enc[4] ^ 
        y_nr_enc[11] ^ 
0; ///1



wire y_nr_47_1;
assign y_nr_47_1 = 
        y_nr_enc[13] ^ 
        y_nr_enc[24] ^ 
        y_nr_enc[36] ^ 
0; ///1



wire y_nr_47_2;
assign y_nr_47_2 = 
        y_nr_enc[43] ^ 
0; ///1



    assign y_nr_p47 = 
y_nr_47_0 ^ 
y_nr_47_1 ^ 
y_nr_47_2 ^ 
0; ///3



wire y_nr_48_0;
assign y_nr_48_0 = 
        y_nr_enc[3] ^ 
        y_nr_enc[14] ^ 
        y_nr_enc[17] ^ 
0; ///1



wire y_nr_48_1;
assign y_nr_48_1 = 
        y_nr_enc[21] ^ 
        y_nr_enc[26] ^ 
        y_nr_enc[28] ^ 
0; ///1



wire y_nr_48_2;
assign y_nr_48_2 = 
        y_nr_enc[32] ^ 
        y_nr_enc[36] ^ 
        y_nr_enc[44] ^ 
0; ///1



    assign y_nr_p48 = 
y_nr_48_0 ^ 
y_nr_48_1 ^ 
y_nr_48_2 ^ 
0; ///3



wire y_nr_49_0;
assign y_nr_49_0 = 
        y_nr_enc[0] ^ 
        y_nr_enc[15] ^ 
        y_nr_enc[18] ^ 
0; ///1



wire y_nr_49_1;
assign y_nr_49_1 = 
        y_nr_enc[22] ^ 
        y_nr_enc[27] ^ 
        y_nr_enc[29] ^ 
0; ///1



wire y_nr_49_2;
assign y_nr_49_2 = 
        y_nr_enc[33] ^ 
        y_nr_enc[37] ^ 
        y_nr_enc[45] ^ 
0; ///1



    assign y_nr_p49 = 
y_nr_49_0 ^ 
y_nr_49_1 ^ 
y_nr_49_2 ^ 
0; ///3



wire y_nr_50_0;
assign y_nr_50_0 = 
        y_nr_enc[1] ^ 
        y_nr_enc[12] ^ 
        y_nr_enc[19] ^ 
0; ///1



wire y_nr_50_1;
assign y_nr_50_1 = 
        y_nr_enc[23] ^ 
        y_nr_enc[24] ^ 
        y_nr_enc[30] ^ 
0; ///1



wire y_nr_50_2;
assign y_nr_50_2 = 
        y_nr_enc[34] ^ 
        y_nr_enc[38] ^ 
        y_nr_enc[46] ^ 
0; ///1



    assign y_nr_p50 = 
y_nr_50_0 ^ 
y_nr_50_1 ^ 
y_nr_50_2 ^ 
0; ///3



wire y_nr_51_0;
assign y_nr_51_0 = 
        y_nr_enc[2] ^ 
        y_nr_enc[13] ^ 
        y_nr_enc[16] ^ 
0; ///1



wire y_nr_51_1;
assign y_nr_51_1 = 
        y_nr_enc[20] ^ 
        y_nr_enc[25] ^ 
        y_nr_enc[31] ^ 
0; ///1



wire y_nr_51_2;
assign y_nr_51_2 = 
        y_nr_enc[35] ^ 
        y_nr_enc[39] ^ 
        y_nr_enc[47] ^ 
0; ///1



    assign y_nr_p51 = 
y_nr_51_0 ^ 
y_nr_51_1 ^ 
y_nr_51_2 ^ 
0; ///3



wire y_nr_52_0;
assign y_nr_52_0 = 
        y_nr_enc[4] ^ 
        y_nr_enc[10] ^ 
        y_nr_enc[18] ^ 
0; ///1



wire y_nr_52_1;
assign y_nr_52_1 = 
        y_nr_enc[20] ^ 
        y_nr_enc[25] ^ 
        y_nr_enc[30] ^ 
0; ///1



wire y_nr_52_2;
assign y_nr_52_2 = 
        y_nr_enc[34] ^ 
        y_nr_enc[36] ^ 
        y_nr_enc[40] ^ 
0; ///1



    assign y_nr_p52 = 
y_nr_52_0 ^ 
y_nr_52_1 ^ 
y_nr_52_2 ^ 
0; ///3



wire y_nr_53_0;
assign y_nr_53_0 = 
        y_nr_enc[5] ^ 
        y_nr_enc[11] ^ 
        y_nr_enc[19] ^ 
0; ///1



wire y_nr_53_1;
assign y_nr_53_1 = 
        y_nr_enc[21] ^ 
        y_nr_enc[26] ^ 
        y_nr_enc[31] ^ 
0; ///1



wire y_nr_53_2;
assign y_nr_53_2 = 
        y_nr_enc[35] ^ 
        y_nr_enc[37] ^ 
        y_nr_enc[41] ^ 
0; ///1



    assign y_nr_p53 = 
y_nr_53_0 ^ 
y_nr_53_1 ^ 
y_nr_53_2 ^ 
0; ///3



wire y_nr_54_0;
assign y_nr_54_0 = 
        y_nr_enc[6] ^ 
        y_nr_enc[8] ^ 
        y_nr_enc[16] ^ 
0; ///1



wire y_nr_54_1;
assign y_nr_54_1 = 
        y_nr_enc[22] ^ 
        y_nr_enc[27] ^ 
        y_nr_enc[28] ^ 
0; ///1



wire y_nr_54_2;
assign y_nr_54_2 = 
        y_nr_enc[32] ^ 
        y_nr_enc[38] ^ 
        y_nr_enc[42] ^ 
0; ///1



    assign y_nr_p54 = 
y_nr_54_0 ^ 
y_nr_54_1 ^ 
y_nr_54_2 ^ 
0; ///3



wire y_nr_55_0;
assign y_nr_55_0 = 
        y_nr_enc[7] ^ 
        y_nr_enc[9] ^ 
        y_nr_enc[17] ^ 
0; ///1



wire y_nr_55_1;
assign y_nr_55_1 = 
        y_nr_enc[23] ^ 
        y_nr_enc[24] ^ 
        y_nr_enc[29] ^ 
0; ///1



wire y_nr_55_2;
assign y_nr_55_2 = 
        y_nr_enc[33] ^ 
        y_nr_enc[39] ^ 
        y_nr_enc[43] ^ 
0; ///1



    assign y_nr_p55 = 
y_nr_55_0 ^ 
y_nr_55_1 ^ 
y_nr_55_2 ^ 
0; ///3



wire y_nr_56_0;
assign y_nr_56_0 = 
        y_nr_enc[3] ^ 
        y_nr_enc[6] ^ 
        y_nr_enc[47] ^ 
0; ///1



    assign y_nr_p56 = 
y_nr_56_0 ^ 
0; ///3



wire y_nr_57_0;
assign y_nr_57_0 = 
        y_nr_enc[0] ^ 
        y_nr_enc[7] ^ 
        y_nr_enc[44] ^ 
0; ///1



    assign y_nr_p57 = 
y_nr_57_0 ^ 
0; ///3



wire y_nr_58_0;
assign y_nr_58_0 = 
        y_nr_enc[1] ^ 
        y_nr_enc[4] ^ 
        y_nr_enc[45] ^ 
0; ///1



    assign y_nr_p58 = 
y_nr_58_0 ^ 
0; ///3



wire y_nr_59_0;
assign y_nr_59_0 = 
        y_nr_enc[2] ^ 
        y_nr_enc[5] ^ 
        y_nr_enc[46] ^ 
0; ///1



    assign y_nr_p59 = 
y_nr_59_0 ^ 
0; ///3



wire y_nr_60_0;
assign y_nr_60_0 = 
        y_nr_enc[3] ^ 
        y_nr_enc[5] ^ 
        y_nr_enc[22] ^ 
0; ///1



wire y_nr_60_1;
assign y_nr_60_1 = 
        y_nr_enc[31] ^ 
        y_nr_enc[47] ^ 
0; ///1



    assign y_nr_p60 = 
y_nr_60_0 ^ 
y_nr_60_1 ^ 
0; ///3



wire y_nr_61_0;
assign y_nr_61_0 = 
        y_nr_enc[0] ^ 
        y_nr_enc[6] ^ 
        y_nr_enc[23] ^ 
0; ///1



wire y_nr_61_1;
assign y_nr_61_1 = 
        y_nr_enc[28] ^ 
        y_nr_enc[44] ^ 
0; ///1



    assign y_nr_p61 = 
y_nr_61_0 ^ 
y_nr_61_1 ^ 
0; ///3



wire y_nr_62_0;
assign y_nr_62_0 = 
        y_nr_enc[1] ^ 
        y_nr_enc[7] ^ 
        y_nr_enc[20] ^ 
0; ///1



wire y_nr_62_1;
assign y_nr_62_1 = 
        y_nr_enc[29] ^ 
        y_nr_enc[45] ^ 
0; ///1



    assign y_nr_p62 = 
y_nr_62_0 ^ 
y_nr_62_1 ^ 
0; ///3



wire y_nr_63_0;
assign y_nr_63_0 = 
        y_nr_enc[2] ^ 
        y_nr_enc[4] ^ 
        y_nr_enc[21] ^ 
0; ///1



wire y_nr_63_1;
assign y_nr_63_1 = 
        y_nr_enc[30] ^ 
        y_nr_enc[46] ^ 
0; ///1



    assign y_nr_p63 = 
y_nr_63_0 ^ 
y_nr_63_1 ^ 
0; ///3



wire y_nr_64_0;
assign y_nr_64_0 = 
        y_nr_enc[3] ^ 
        y_nr_enc[20] ^ 
        y_nr_enc[29] ^ 
0; ///1



wire y_nr_64_1;
assign y_nr_64_1 = 
        y_nr_enc[36] ^ 
        y_nr_enc[46] ^ 
0; ///1



    assign y_nr_p64 = 
y_nr_64_0 ^ 
y_nr_64_1 ^ 
0; ///3



wire y_nr_65_0;
assign y_nr_65_0 = 
        y_nr_enc[0] ^ 
        y_nr_enc[21] ^ 
        y_nr_enc[30] ^ 
0; ///1



wire y_nr_65_1;
assign y_nr_65_1 = 
        y_nr_enc[37] ^ 
        y_nr_enc[47] ^ 
0; ///1



    assign y_nr_p65 = 
y_nr_65_0 ^ 
y_nr_65_1 ^ 
0; ///3



wire y_nr_66_0;
assign y_nr_66_0 = 
        y_nr_enc[1] ^ 
        y_nr_enc[22] ^ 
        y_nr_enc[31] ^ 
0; ///1



wire y_nr_66_1;
assign y_nr_66_1 = 
        y_nr_enc[38] ^ 
        y_nr_enc[44] ^ 
0; ///1



    assign y_nr_p66 = 
y_nr_66_0 ^ 
y_nr_66_1 ^ 
0; ///3



wire y_nr_67_0;
assign y_nr_67_0 = 
        y_nr_enc[2] ^ 
        y_nr_enc[23] ^ 
        y_nr_enc[28] ^ 
0; ///1



wire y_nr_67_1;
assign y_nr_67_1 = 
        y_nr_enc[39] ^ 
        y_nr_enc[45] ^ 
0; ///1



    assign y_nr_p67 = 
y_nr_67_0 ^ 
y_nr_67_1 ^ 
0; ///3



wire y_nr_68_0;
assign y_nr_68_0 = 
        y_nr_enc[5] ^ 
        y_nr_enc[23] ^ 
        y_nr_enc[28] ^ 
0; ///1



wire y_nr_68_1;
assign y_nr_68_1 = 
        y_nr_enc[47] ^ 
        y_nr_enc[52] ^ 
0; ///1



    assign y_nr_p68 = 
y_nr_68_0 ^ 
y_nr_68_1 ^ 
0; ///3



wire y_nr_69_0;
assign y_nr_69_0 = 
        y_nr_enc[6] ^ 
        y_nr_enc[20] ^ 
        y_nr_enc[29] ^ 
0; ///1



wire y_nr_69_1;
assign y_nr_69_1 = 
        y_nr_enc[44] ^ 
        y_nr_enc[53] ^ 
0; ///1



    assign y_nr_p69 = 
y_nr_69_0 ^ 
y_nr_69_1 ^ 
0; ///3



wire y_nr_70_0;
assign y_nr_70_0 = 
        y_nr_enc[7] ^ 
        y_nr_enc[21] ^ 
        y_nr_enc[30] ^ 
0; ///1



wire y_nr_70_1;
assign y_nr_70_1 = 
        y_nr_enc[45] ^ 
        y_nr_enc[54] ^ 
0; ///1



    assign y_nr_p70 = 
y_nr_70_0 ^ 
y_nr_70_1 ^ 
0; ///3



wire y_nr_71_0;
assign y_nr_71_0 = 
        y_nr_enc[4] ^ 
        y_nr_enc[22] ^ 
        y_nr_enc[31] ^ 
0; ///1



wire y_nr_71_1;
assign y_nr_71_1 = 
        y_nr_enc[46] ^ 
        y_nr_enc[55] ^ 
0; ///1



    assign y_nr_p71 = 
y_nr_71_0 ^ 
y_nr_71_1 ^ 
0; ///3



wire y_nr_72_0;
assign y_nr_72_0 = 
        y_nr_enc[2] ^ 
        y_nr_enc[6] ^ 
        y_nr_enc[50] ^ 
0; ///1



    assign y_nr_p72 = 
y_nr_72_0 ^ 
0; ///3



wire y_nr_73_0;
assign y_nr_73_0 = 
        y_nr_enc[3] ^ 
        y_nr_enc[7] ^ 
        y_nr_enc[51] ^ 
0; ///1



    assign y_nr_p73 = 
y_nr_73_0 ^ 
0; ///3



wire y_nr_74_0;
assign y_nr_74_0 = 
        y_nr_enc[0] ^ 
        y_nr_enc[4] ^ 
        y_nr_enc[48] ^ 
0; ///1



    assign y_nr_p74 = 
y_nr_74_0 ^ 
0; ///3



wire y_nr_75_0;
assign y_nr_75_0 = 
        y_nr_enc[1] ^ 
        y_nr_enc[5] ^ 
        y_nr_enc[49] ^ 
0; ///1



    assign y_nr_p75 = 
y_nr_75_0 ^ 
0; ///3



wire y_nr_76_0;
assign y_nr_76_0 = 
        y_nr_enc[7] ^ 
        y_nr_enc[33] ^ 
        y_nr_enc[41] ^ 
0; ///1



wire y_nr_76_1;
assign y_nr_76_1 = 
        y_nr_enc[47] ^ 
0; ///1



    assign y_nr_p76 = 
y_nr_76_0 ^ 
y_nr_76_1 ^ 
0; ///3



wire y_nr_77_0;
assign y_nr_77_0 = 
        y_nr_enc[4] ^ 
        y_nr_enc[34] ^ 
        y_nr_enc[42] ^ 
0; ///1



wire y_nr_77_1;
assign y_nr_77_1 = 
        y_nr_enc[44] ^ 
0; ///1



    assign y_nr_p77 = 
y_nr_77_0 ^ 
y_nr_77_1 ^ 
0; ///3



wire y_nr_78_0;
assign y_nr_78_0 = 
        y_nr_enc[5] ^ 
        y_nr_enc[35] ^ 
        y_nr_enc[43] ^ 
0; ///1



wire y_nr_78_1;
assign y_nr_78_1 = 
        y_nr_enc[45] ^ 
0; ///1



    assign y_nr_p78 = 
y_nr_78_0 ^ 
y_nr_78_1 ^ 
0; ///3



wire y_nr_79_0;
assign y_nr_79_0 = 
        y_nr_enc[6] ^ 
        y_nr_enc[32] ^ 
        y_nr_enc[40] ^ 
0; ///1



wire y_nr_79_1;
assign y_nr_79_1 = 
        y_nr_enc[46] ^ 
0; ///1



    assign y_nr_p79 = 
y_nr_79_0 ^ 
y_nr_79_1 ^ 
0; ///3



wire y_nr_80_0;
assign y_nr_80_0 = 
        y_nr_enc[3] ^ 
        y_nr_enc[5] ^ 
        y_nr_enc[24] ^ 
0; ///1



wire y_nr_80_1;
assign y_nr_80_1 = 
        y_nr_enc[29] ^ 
0; ///1



    assign y_nr_p80 = 
y_nr_80_0 ^ 
y_nr_80_1 ^ 
0; ///3



wire y_nr_81_0;
assign y_nr_81_0 = 
        y_nr_enc[0] ^ 
        y_nr_enc[6] ^ 
        y_nr_enc[25] ^ 
0; ///1



wire y_nr_81_1;
assign y_nr_81_1 = 
        y_nr_enc[30] ^ 
0; ///1



    assign y_nr_p81 = 
y_nr_81_0 ^ 
y_nr_81_1 ^ 
0; ///3



wire y_nr_82_0;
assign y_nr_82_0 = 
        y_nr_enc[1] ^ 
        y_nr_enc[7] ^ 
        y_nr_enc[26] ^ 
0; ///1



wire y_nr_82_1;
assign y_nr_82_1 = 
        y_nr_enc[31] ^ 
0; ///1



    assign y_nr_p82 = 
y_nr_82_0 ^ 
y_nr_82_1 ^ 
0; ///3



wire y_nr_83_0;
assign y_nr_83_0 = 
        y_nr_enc[2] ^ 
        y_nr_enc[4] ^ 
        y_nr_enc[27] ^ 
0; ///1



wire y_nr_83_1;
assign y_nr_83_1 = 
        y_nr_enc[28] ^ 
0; ///1



    assign y_nr_p83 = 
y_nr_83_0 ^ 
y_nr_83_1 ^ 
0; ///3



wire y_nr_84_0;
assign y_nr_84_0 = 
        y_nr_enc[3] ^ 
        y_nr_enc[28] ^ 
        y_nr_enc[38] ^ 
0; ///1



wire y_nr_84_1;
assign y_nr_84_1 = 
        y_nr_enc[52] ^ 
0; ///1



    assign y_nr_p84 = 
y_nr_84_0 ^ 
y_nr_84_1 ^ 
0; ///3



wire y_nr_85_0;
assign y_nr_85_0 = 
        y_nr_enc[0] ^ 
        y_nr_enc[29] ^ 
        y_nr_enc[39] ^ 
0; ///1



wire y_nr_85_1;
assign y_nr_85_1 = 
        y_nr_enc[53] ^ 
0; ///1



    assign y_nr_p85 = 
y_nr_85_0 ^ 
y_nr_85_1 ^ 
0; ///3



wire y_nr_86_0;
assign y_nr_86_0 = 
        y_nr_enc[1] ^ 
        y_nr_enc[30] ^ 
        y_nr_enc[36] ^ 
0; ///1



wire y_nr_86_1;
assign y_nr_86_1 = 
        y_nr_enc[54] ^ 
0; ///1



    assign y_nr_p86 = 
y_nr_86_0 ^ 
y_nr_86_1 ^ 
0; ///3



wire y_nr_87_0;
assign y_nr_87_0 = 
        y_nr_enc[2] ^ 
        y_nr_enc[31] ^ 
        y_nr_enc[37] ^ 
0; ///1



wire y_nr_87_1;
assign y_nr_87_1 = 
        y_nr_enc[55] ^ 
0; ///1



    assign y_nr_p87 = 
y_nr_87_0 ^ 
y_nr_87_1 ^ 
0; ///3



wire y_nr_88_0;
assign y_nr_88_0 = 
        y_nr_enc[7] ^ 
        y_nr_enc[15] ^ 
        y_nr_enc[46] ^ 
0; ///1



    assign y_nr_p88 = 
y_nr_88_0 ^ 
0; ///3



wire y_nr_89_0;
assign y_nr_89_0 = 
        y_nr_enc[4] ^ 
        y_nr_enc[12] ^ 
        y_nr_enc[47] ^ 
0; ///1



    assign y_nr_p89 = 
y_nr_89_0 ^ 
0; ///3



wire y_nr_90_0;
assign y_nr_90_0 = 
        y_nr_enc[5] ^ 
        y_nr_enc[13] ^ 
        y_nr_enc[44] ^ 
0; ///1



    assign y_nr_p90 = 
y_nr_90_0 ^ 
0; ///3



wire y_nr_91_0;
assign y_nr_91_0 = 
        y_nr_enc[6] ^ 
        y_nr_enc[14] ^ 
        y_nr_enc[45] ^ 
0; ///1



    assign y_nr_p91 = 
y_nr_91_0 ^ 
0; ///3



wire y_nr_92_0;
assign y_nr_92_0 = 
        y_nr_enc[3] ^ 
        y_nr_enc[6] ^ 
        y_nr_enc[34] ^ 
0; ///1



wire y_nr_92_1;
assign y_nr_92_1 = 
        y_nr_enc[54] ^ 
0; ///1



    assign y_nr_p92 = 
y_nr_92_0 ^ 
y_nr_92_1 ^ 
0; ///3



wire y_nr_93_0;
assign y_nr_93_0 = 
        y_nr_enc[0] ^ 
        y_nr_enc[7] ^ 
        y_nr_enc[35] ^ 
0; ///1



wire y_nr_93_1;
assign y_nr_93_1 = 
        y_nr_enc[55] ^ 
0; ///1



    assign y_nr_p93 = 
y_nr_93_0 ^ 
y_nr_93_1 ^ 
0; ///3



wire y_nr_94_0;
assign y_nr_94_0 = 
        y_nr_enc[1] ^ 
        y_nr_enc[4] ^ 
        y_nr_enc[32] ^ 
0; ///1



wire y_nr_94_1;
assign y_nr_94_1 = 
        y_nr_enc[52] ^ 
0; ///1



    assign y_nr_p94 = 
y_nr_94_0 ^ 
y_nr_94_1 ^ 
0; ///3



wire y_nr_95_0;
assign y_nr_95_0 = 
        y_nr_enc[2] ^ 
        y_nr_enc[5] ^ 
        y_nr_enc[33] ^ 
0; ///1



wire y_nr_95_1;
assign y_nr_95_1 = 
        y_nr_enc[53] ^ 
0; ///1



    assign y_nr_p95 = 
y_nr_95_0 ^ 
y_nr_95_1 ^ 
0; ///3



wire y_nr_96_0;
assign y_nr_96_0 = 
        y_nr_enc[7] ^ 
        y_nr_enc[25] ^ 
        y_nr_enc[47] ^ 
0; ///1



wire y_nr_96_1;
assign y_nr_96_1 = 
        y_nr_enc[52] ^ 
0; ///1



    assign y_nr_p96 = 
y_nr_96_0 ^ 
y_nr_96_1 ^ 
0; ///3



wire y_nr_97_0;
assign y_nr_97_0 = 
        y_nr_enc[4] ^ 
        y_nr_enc[26] ^ 
        y_nr_enc[44] ^ 
0; ///1



wire y_nr_97_1;
assign y_nr_97_1 = 
        y_nr_enc[53] ^ 
0; ///1



    assign y_nr_p97 = 
y_nr_97_0 ^ 
y_nr_97_1 ^ 
0; ///3



wire y_nr_98_0;
assign y_nr_98_0 = 
        y_nr_enc[5] ^ 
        y_nr_enc[27] ^ 
        y_nr_enc[45] ^ 
0; ///1



wire y_nr_98_1;
assign y_nr_98_1 = 
        y_nr_enc[54] ^ 
0; ///1



    assign y_nr_p98 = 
y_nr_98_0 ^ 
y_nr_98_1 ^ 
0; ///3



wire y_nr_99_0;
assign y_nr_99_0 = 
        y_nr_enc[6] ^ 
        y_nr_enc[24] ^ 
        y_nr_enc[46] ^ 
0; ///1



wire y_nr_99_1;
assign y_nr_99_1 = 
        y_nr_enc[55] ^ 
0; ///1



    assign y_nr_p99 = 
y_nr_99_0 ^ 
y_nr_99_1 ^ 
0; ///3



wire y_nr_100_0;
assign y_nr_100_0 = 
        y_nr_enc[3] ^ 
        y_nr_enc[43] ^ 
        y_nr_enc[45] ^ 
0; ///1



    assign y_nr_p100 = 
y_nr_100_0 ^ 
0; ///3



wire y_nr_101_0;
assign y_nr_101_0 = 
        y_nr_enc[0] ^ 
        y_nr_enc[40] ^ 
        y_nr_enc[46] ^ 
0; ///1



    assign y_nr_p101 = 
y_nr_101_0 ^ 
0; ///3



wire y_nr_102_0;
assign y_nr_102_0 = 
        y_nr_enc[1] ^ 
        y_nr_enc[41] ^ 
        y_nr_enc[47] ^ 
0; ///1



    assign y_nr_p102 = 
y_nr_102_0 ^ 
0; ///3



wire y_nr_103_0;
assign y_nr_103_0 = 
        y_nr_enc[2] ^ 
        y_nr_enc[42] ^ 
        y_nr_enc[44] ^ 
0; ///1



    assign y_nr_p103 = 
y_nr_103_0 ^ 
0; ///3



wire y_nr_104_0;
assign y_nr_104_0 = 
        y_nr_enc[7] ^ 
        y_nr_enc[38] ^ 
        y_nr_enc[44] ^ 
0; ///1



wire y_nr_104_1;
assign y_nr_104_1 = 
        y_nr_enc[50] ^ 
0; ///1



    assign y_nr_p104 = 
y_nr_104_0 ^ 
y_nr_104_1 ^ 
0; ///3



wire y_nr_105_0;
assign y_nr_105_0 = 
        y_nr_enc[4] ^ 
        y_nr_enc[39] ^ 
        y_nr_enc[45] ^ 
0; ///1



wire y_nr_105_1;
assign y_nr_105_1 = 
        y_nr_enc[51] ^ 
0; ///1



    assign y_nr_p105 = 
y_nr_105_0 ^ 
y_nr_105_1 ^ 
0; ///3



wire y_nr_106_0;
assign y_nr_106_0 = 
        y_nr_enc[5] ^ 
        y_nr_enc[36] ^ 
        y_nr_enc[46] ^ 
0; ///1



wire y_nr_106_1;
assign y_nr_106_1 = 
        y_nr_enc[48] ^ 
0; ///1



    assign y_nr_p106 = 
y_nr_106_0 ^ 
y_nr_106_1 ^ 
0; ///3



wire y_nr_107_0;
assign y_nr_107_0 = 
        y_nr_enc[6] ^ 
        y_nr_enc[37] ^ 
        y_nr_enc[47] ^ 
0; ///1



wire y_nr_107_1;
assign y_nr_107_1 = 
        y_nr_enc[49] ^ 
0; ///1



    assign y_nr_p107 = 
y_nr_107_0 ^ 
y_nr_107_1 ^ 
0; ///3



wire y_nr_108_0;
assign y_nr_108_0 = 
        y_nr_enc[6] ^ 
        y_nr_enc[20] ^ 
        y_nr_enc[46] ^ 
0; ///1



wire y_nr_108_1;
assign y_nr_108_1 = 
        y_nr_enc[48] ^ 
0; ///1



    assign y_nr_p108 = 
y_nr_108_0 ^ 
y_nr_108_1 ^ 
0; ///3



wire y_nr_109_0;
assign y_nr_109_0 = 
        y_nr_enc[7] ^ 
        y_nr_enc[21] ^ 
        y_nr_enc[47] ^ 
0; ///1



wire y_nr_109_1;
assign y_nr_109_1 = 
        y_nr_enc[49] ^ 
0; ///1



    assign y_nr_p109 = 
y_nr_109_0 ^ 
y_nr_109_1 ^ 
0; ///3



wire y_nr_110_0;
assign y_nr_110_0 = 
        y_nr_enc[4] ^ 
        y_nr_enc[22] ^ 
        y_nr_enc[44] ^ 
0; ///1



wire y_nr_110_1;
assign y_nr_110_1 = 
        y_nr_enc[50] ^ 
0; ///1



    assign y_nr_p110 = 
y_nr_110_0 ^ 
y_nr_110_1 ^ 
0; ///3



wire y_nr_111_0;
assign y_nr_111_0 = 
        y_nr_enc[5] ^ 
        y_nr_enc[23] ^ 
        y_nr_enc[45] ^ 
0; ///1



wire y_nr_111_1;
assign y_nr_111_1 = 
        y_nr_enc[51] ^ 
0; ///1



    assign y_nr_p111 = 
y_nr_111_0 ^ 
y_nr_111_1 ^ 
0; ///3



wire y_nr_112_0;
assign y_nr_112_0 = 
        y_nr_enc[0] ^ 
        y_nr_enc[26] ^ 
        y_nr_enc[30] ^ 
0; ///1



    assign y_nr_p112 = 
y_nr_112_0 ^ 
0; ///3



wire y_nr_113_0;
assign y_nr_113_0 = 
        y_nr_enc[1] ^ 
        y_nr_enc[27] ^ 
        y_nr_enc[31] ^ 
0; ///1



    assign y_nr_p113 = 
y_nr_113_0 ^ 
0; ///3



wire y_nr_114_0;
assign y_nr_114_0 = 
        y_nr_enc[2] ^ 
        y_nr_enc[24] ^ 
        y_nr_enc[28] ^ 
0; ///1



    assign y_nr_p114 = 
y_nr_114_0 ^ 
0; ///3



wire y_nr_115_0;
assign y_nr_115_0 = 
        y_nr_enc[3] ^ 
        y_nr_enc[25] ^ 
        y_nr_enc[29] ^ 
0; ///1



    assign y_nr_p115 = 
y_nr_115_0 ^ 
0; ///3



wire y_nr_116_0;
assign y_nr_116_0 = 
        y_nr_enc[3] ^ 
        y_nr_enc[4] ^ 
        y_nr_enc[41] ^ 
0; ///1



    assign y_nr_p116 = 
y_nr_116_0 ^ 
0; ///3



wire y_nr_117_0;
assign y_nr_117_0 = 
        y_nr_enc[0] ^ 
        y_nr_enc[5] ^ 
        y_nr_enc[42] ^ 
0; ///1



    assign y_nr_p117 = 
y_nr_117_0 ^ 
0; ///3



wire y_nr_118_0;
assign y_nr_118_0 = 
        y_nr_enc[1] ^ 
        y_nr_enc[6] ^ 
        y_nr_enc[43] ^ 
0; ///1



    assign y_nr_p118 = 
y_nr_118_0 ^ 
0; ///3



wire y_nr_119_0;
assign y_nr_119_0 = 
        y_nr_enc[2] ^ 
        y_nr_enc[7] ^ 
        y_nr_enc[40] ^ 
0; ///1



    assign y_nr_p119 = 
y_nr_119_0 ^ 
0; ///3



wire y_nr_120_0;
assign y_nr_120_0 = 
        y_nr_enc[6] ^ 
        y_nr_enc[17] ^ 
        y_nr_enc[45] ^ 
0; ///1



    assign y_nr_p120 = 
y_nr_120_0 ^ 
0; ///3



wire y_nr_121_0;
assign y_nr_121_0 = 
        y_nr_enc[7] ^ 
        y_nr_enc[18] ^ 
        y_nr_enc[46] ^ 
0; ///1



    assign y_nr_p121 = 
y_nr_121_0 ^ 
0; ///3



wire y_nr_122_0;
assign y_nr_122_0 = 
        y_nr_enc[4] ^ 
        y_nr_enc[19] ^ 
        y_nr_enc[47] ^ 
0; ///1



    assign y_nr_p122 = 
y_nr_122_0 ^ 
0; ///3



wire y_nr_123_0;
assign y_nr_123_0 = 
        y_nr_enc[5] ^ 
        y_nr_enc[16] ^ 
        y_nr_enc[44] ^ 
0; ///1



    assign y_nr_p123 = 
y_nr_123_0 ^ 
0; ///3



wire y_nr_124_0;
assign y_nr_124_0 = 
        y_nr_enc[0] ^ 
        y_nr_enc[34] ^ 
        y_nr_enc[54] ^ 
0; ///1



    assign y_nr_p124 = 
y_nr_124_0 ^ 
0; ///3



wire y_nr_125_0;
assign y_nr_125_0 = 
        y_nr_enc[1] ^ 
        y_nr_enc[35] ^ 
        y_nr_enc[55] ^ 
0; ///1



    assign y_nr_p125 = 
y_nr_125_0 ^ 
0; ///3



wire y_nr_126_0;
assign y_nr_126_0 = 
        y_nr_enc[2] ^ 
        y_nr_enc[32] ^ 
        y_nr_enc[52] ^ 
0; ///1



    assign y_nr_p126 = 
y_nr_126_0 ^ 
0; ///3



wire y_nr_127_0;
assign y_nr_127_0 = 
        y_nr_enc[3] ^ 
        y_nr_enc[33] ^ 
        y_nr_enc[53] ^ 
0; ///1



    assign y_nr_p127 = 
y_nr_127_0 ^ 
0; ///3



wire y_nr_128_0;
assign y_nr_128_0 = 
        y_nr_enc[6] ^ 
        y_nr_enc[11] ^ 
0; ///1



    assign y_nr_p128 = 
y_nr_128_0 ^ 
0; ///3



wire y_nr_129_0;
assign y_nr_129_0 = 
        y_nr_enc[7] ^ 
        y_nr_enc[8] ^ 
0; ///1



    assign y_nr_p129 = 
y_nr_129_0 ^ 
0; ///3



wire y_nr_130_0;
assign y_nr_130_0 = 
        y_nr_enc[4] ^ 
        y_nr_enc[9] ^ 
0; ///1



    assign y_nr_p130 = 
y_nr_130_0 ^ 
0; ///3



wire y_nr_131_0;
assign y_nr_131_0 = 
        y_nr_enc[5] ^ 
        y_nr_enc[10] ^ 
0; ///1



    assign y_nr_p131 = 
y_nr_131_0 ^ 
0; ///3



wire y_nr_132_0;
assign y_nr_132_0 = 
        y_nr_enc[3] ^ 
        y_nr_enc[15] ^ 
        y_nr_enc[22] ^ 
0; ///1



    assign y_nr_p132 = 
y_nr_132_0 ^ 
0; ///3



wire y_nr_133_0;
assign y_nr_133_0 = 
        y_nr_enc[0] ^ 
        y_nr_enc[12] ^ 
        y_nr_enc[23] ^ 
0; ///1



    assign y_nr_p133 = 
y_nr_133_0 ^ 
0; ///3



wire y_nr_134_0;
assign y_nr_134_0 = 
        y_nr_enc[1] ^ 
        y_nr_enc[13] ^ 
        y_nr_enc[20] ^ 
0; ///1



    assign y_nr_p134 = 
y_nr_134_0 ^ 
0; ///3



wire y_nr_135_0;
assign y_nr_135_0 = 
        y_nr_enc[2] ^ 
        y_nr_enc[14] ^ 
        y_nr_enc[21] ^ 
0; ///1



    assign y_nr_p135 = 
y_nr_135_0 ^ 
0; ///3



wire y_nr_136_0;
assign y_nr_136_0 = 
        y_nr_enc[6] ^ 
        y_nr_enc[11] ^ 
        y_nr_enc[36] ^ 
0; ///1



    assign y_nr_p136 = 
y_nr_136_0 ^ 
0; ///3



wire y_nr_137_0;
assign y_nr_137_0 = 
        y_nr_enc[7] ^ 
        y_nr_enc[8] ^ 
        y_nr_enc[37] ^ 
0; ///1



    assign y_nr_p137 = 
y_nr_137_0 ^ 
0; ///3



wire y_nr_138_0;
assign y_nr_138_0 = 
        y_nr_enc[4] ^ 
        y_nr_enc[9] ^ 
        y_nr_enc[38] ^ 
0; ///1



    assign y_nr_p138 = 
y_nr_138_0 ^ 
0; ///3



wire y_nr_139_0;
assign y_nr_139_0 = 
        y_nr_enc[5] ^ 
        y_nr_enc[10] ^ 
        y_nr_enc[39] ^ 
0; ///1



    assign y_nr_p139 = 
y_nr_139_0 ^ 
0; ///3



wire y_nr_140_0;
assign y_nr_140_0 = 
        y_nr_enc[0] ^ 
        y_nr_enc[20] ^ 
0; ///1



    assign y_nr_p140 = 
y_nr_140_0 ^ 
0; ///3



wire y_nr_141_0;
assign y_nr_141_0 = 
        y_nr_enc[1] ^ 
        y_nr_enc[21] ^ 
0; ///1



    assign y_nr_p141 = 
y_nr_141_0 ^ 
0; ///3



wire y_nr_142_0;
assign y_nr_142_0 = 
        y_nr_enc[2] ^ 
        y_nr_enc[22] ^ 
0; ///1



    assign y_nr_p142 = 
y_nr_142_0 ^ 
0; ///3



wire y_nr_143_0;
assign y_nr_143_0 = 
        y_nr_enc[3] ^ 
        y_nr_enc[23] ^ 
0; ///1



    assign y_nr_p143 = 
y_nr_143_0 ^ 
0; ///3



wire y_nr_144_0;
assign y_nr_144_0 = 
        y_nr_enc[9] ^ 
        y_nr_enc[31] ^ 
        y_nr_enc[48] ^ 
0; ///1



wire y_nr_144_1;
assign y_nr_144_1 = 
        y_nr_enc[54] ^ 
0; ///1



    assign y_nr_p144 = 
y_nr_144_0 ^ 
y_nr_144_1 ^ 
0; ///3



wire y_nr_145_0;
assign y_nr_145_0 = 
        y_nr_enc[10] ^ 
        y_nr_enc[28] ^ 
        y_nr_enc[49] ^ 
0; ///1



wire y_nr_145_1;
assign y_nr_145_1 = 
        y_nr_enc[55] ^ 
0; ///1



    assign y_nr_p145 = 
y_nr_145_0 ^ 
y_nr_145_1 ^ 
0; ///3



wire y_nr_146_0;
assign y_nr_146_0 = 
        y_nr_enc[11] ^ 
        y_nr_enc[29] ^ 
        y_nr_enc[50] ^ 
0; ///1



wire y_nr_146_1;
assign y_nr_146_1 = 
        y_nr_enc[52] ^ 
0; ///1



    assign y_nr_p146 = 
y_nr_146_0 ^ 
y_nr_146_1 ^ 
0; ///3



wire y_nr_147_0;
assign y_nr_147_0 = 
        y_nr_enc[8] ^ 
        y_nr_enc[30] ^ 
        y_nr_enc[51] ^ 
0; ///1



wire y_nr_147_1;
assign y_nr_147_1 = 
        y_nr_enc[53] ^ 
0; ///1



    assign y_nr_p147 = 
y_nr_147_0 ^ 
y_nr_147_1 ^ 
0; ///3



wire y_nr_148_0;
assign y_nr_148_0 = 
        y_nr_enc[0] ^ 
        y_nr_enc[27] ^ 
0; ///1



    assign y_nr_p148 = 
y_nr_148_0 ^ 
0; ///3



wire y_nr_149_0;
assign y_nr_149_0 = 
        y_nr_enc[1] ^ 
        y_nr_enc[24] ^ 
0; ///1



    assign y_nr_p149 = 
y_nr_149_0 ^ 
0; ///3



wire y_nr_150_0;
assign y_nr_150_0 = 
        y_nr_enc[2] ^ 
        y_nr_enc[25] ^ 
0; ///1



    assign y_nr_p150 = 
y_nr_150_0 ^ 
0; ///3



wire y_nr_151_0;
assign y_nr_151_0 = 
        y_nr_enc[3] ^ 
        y_nr_enc[26] ^ 
0; ///1



    assign y_nr_p151 = 
y_nr_151_0 ^ 
0; ///3



wire y_nr_152_0;
assign y_nr_152_0 = 
        y_nr_enc[6] ^ 
        y_nr_enc[9] ^ 
        y_nr_enc[23] ^ 
0; ///1



    assign y_nr_p152 = 
y_nr_152_0 ^ 
0; ///3



wire y_nr_153_0;
assign y_nr_153_0 = 
        y_nr_enc[7] ^ 
        y_nr_enc[10] ^ 
        y_nr_enc[20] ^ 
0; ///1



    assign y_nr_p153 = 
y_nr_153_0 ^ 
0; ///3



wire y_nr_154_0;
assign y_nr_154_0 = 
        y_nr_enc[4] ^ 
        y_nr_enc[11] ^ 
        y_nr_enc[21] ^ 
0; ///1



    assign y_nr_p154 = 
y_nr_154_0 ^ 
0; ///3



wire y_nr_155_0;
assign y_nr_155_0 = 
        y_nr_enc[5] ^ 
        y_nr_enc[8] ^ 
        y_nr_enc[22] ^ 
0; ///1



    assign y_nr_p155 = 
y_nr_155_0 ^ 
0; ///3



wire y_nr_156_0;
assign y_nr_156_0 = 
        y_nr_enc[2] ^ 
        y_nr_enc[16] ^ 
0; ///1



    assign y_nr_p156 = 
y_nr_156_0 ^ 
0; ///3



wire y_nr_157_0;
assign y_nr_157_0 = 
        y_nr_enc[3] ^ 
        y_nr_enc[17] ^ 
0; ///1



    assign y_nr_p157 = 
y_nr_157_0 ^ 
0; ///3



wire y_nr_158_0;
assign y_nr_158_0 = 
        y_nr_enc[0] ^ 
        y_nr_enc[18] ^ 
0; ///1



    assign y_nr_p158 = 
y_nr_158_0 ^ 
0; ///3



wire y_nr_159_0;
assign y_nr_159_0 = 
        y_nr_enc[1] ^ 
        y_nr_enc[19] ^ 
0; ///1



    assign y_nr_p159 = 
y_nr_159_0 ^ 
0; ///3



wire y_nr_160_0;
assign y_nr_160_0 = 
        y_nr_enc[11] ^ 
        y_nr_enc[20] ^ 
        y_nr_enc[29] ^ 
0; ///1



wire y_nr_160_1;
assign y_nr_160_1 = 
        y_nr_enc[36] ^ 
0; ///1



    assign y_nr_p160 = 
y_nr_160_0 ^ 
y_nr_160_1 ^ 
0; ///3



wire y_nr_161_0;
assign y_nr_161_0 = 
        y_nr_enc[8] ^ 
        y_nr_enc[21] ^ 
        y_nr_enc[30] ^ 
0; ///1



wire y_nr_161_1;
assign y_nr_161_1 = 
        y_nr_enc[37] ^ 
0; ///1



    assign y_nr_p161 = 
y_nr_161_0 ^ 
y_nr_161_1 ^ 
0; ///3



wire y_nr_162_0;
assign y_nr_162_0 = 
        y_nr_enc[9] ^ 
        y_nr_enc[22] ^ 
        y_nr_enc[31] ^ 
0; ///1



wire y_nr_162_1;
assign y_nr_162_1 = 
        y_nr_enc[38] ^ 
0; ///1



    assign y_nr_p162 = 
y_nr_162_0 ^ 
y_nr_162_1 ^ 
0; ///3



wire y_nr_163_0;
assign y_nr_163_0 = 
        y_nr_enc[10] ^ 
        y_nr_enc[23] ^ 
        y_nr_enc[28] ^ 
0; ///1



wire y_nr_163_1;
assign y_nr_163_1 = 
        y_nr_enc[39] ^ 
0; ///1



    assign y_nr_p163 = 
y_nr_163_0 ^ 
y_nr_163_1 ^ 
0; ///3



wire y_nr_164_0;
assign y_nr_164_0 = 
        y_nr_enc[6] ^ 
        y_nr_enc[53] ^ 
0; ///1



    assign y_nr_p164 = 
y_nr_164_0 ^ 
0; ///3



wire y_nr_165_0;
assign y_nr_165_0 = 
        y_nr_enc[7] ^ 
        y_nr_enc[54] ^ 
0; ///1



    assign y_nr_p165 = 
y_nr_165_0 ^ 
0; ///3



wire y_nr_166_0;
assign y_nr_166_0 = 
        y_nr_enc[4] ^ 
        y_nr_enc[55] ^ 
0; ///1



    assign y_nr_p166 = 
y_nr_166_0 ^ 
0; ///3



wire y_nr_167_0;
assign y_nr_167_0 = 
        y_nr_enc[5] ^ 
        y_nr_enc[52] ^ 
0; ///1



    assign y_nr_p167 = 
y_nr_167_0 ^ 
0; ///3



wire y_nr_168_0;
assign y_nr_168_0 = 
        y_nr_enc[2] ^ 
        y_nr_enc[20] ^ 
        y_nr_enc[50] ^ 
0; ///1



    assign y_nr_p168 = 
y_nr_168_0 ^ 
0; ///3



wire y_nr_169_0;
assign y_nr_169_0 = 
        y_nr_enc[3] ^ 
        y_nr_enc[21] ^ 
        y_nr_enc[51] ^ 
0; ///1



    assign y_nr_p169 = 
y_nr_169_0 ^ 
0; ///3



wire y_nr_170_0;
assign y_nr_170_0 = 
        y_nr_enc[0] ^ 
        y_nr_enc[22] ^ 
        y_nr_enc[48] ^ 
0; ///1



    assign y_nr_p170 = 
y_nr_170_0 ^ 
0; ///3



wire y_nr_171_0;
assign y_nr_171_0 = 
        y_nr_enc[1] ^ 
        y_nr_enc[23] ^ 
        y_nr_enc[49] ^ 
0; ///1



    assign y_nr_p171 = 
y_nr_171_0 ^ 
0; ///3



wire y_nr_172_0;
assign y_nr_172_0 = 
        y_nr_enc[8] ^ 
        y_nr_enc[28] ^ 
        y_nr_enc[43] ^ 
0; ///1



    assign y_nr_p172 = 
y_nr_172_0 ^ 
0; ///3



wire y_nr_173_0;
assign y_nr_173_0 = 
        y_nr_enc[9] ^ 
        y_nr_enc[29] ^ 
        y_nr_enc[40] ^ 
0; ///1



    assign y_nr_p173 = 
y_nr_173_0 ^ 
0; ///3



wire y_nr_174_0;
assign y_nr_174_0 = 
        y_nr_enc[10] ^ 
        y_nr_enc[30] ^ 
        y_nr_enc[41] ^ 
0; ///1



    assign y_nr_p174 = 
y_nr_174_0 ^ 
0; ///3



wire y_nr_175_0;
assign y_nr_175_0 = 
        y_nr_enc[11] ^ 
        y_nr_enc[31] ^ 
        y_nr_enc[42] ^ 
0; ///1



    assign y_nr_p175 = 
y_nr_175_0 ^ 
0; ///3



wire y_nr_176_0;
assign y_nr_176_0 = 
        y_nr_enc[3] ^ 
        y_nr_enc[49] ^ 
        y_nr_enc[52] ^ 
0; ///1



    assign y_nr_p176 = 
y_nr_176_0 ^ 
0; ///3



wire y_nr_177_0;
assign y_nr_177_0 = 
        y_nr_enc[0] ^ 
        y_nr_enc[50] ^ 
        y_nr_enc[53] ^ 
0; ///1



    assign y_nr_p177 = 
y_nr_177_0 ^ 
0; ///3



wire y_nr_178_0;
assign y_nr_178_0 = 
        y_nr_enc[1] ^ 
        y_nr_enc[51] ^ 
        y_nr_enc[54] ^ 
0; ///1



    assign y_nr_p178 = 
y_nr_178_0 ^ 
0; ///3



wire y_nr_179_0;
assign y_nr_179_0 = 
        y_nr_enc[2] ^ 
        y_nr_enc[48] ^ 
        y_nr_enc[55] ^ 
0; ///1



    assign y_nr_p179 = 
y_nr_179_0 ^ 
0; ///3



wire y_nr_180_0;
assign y_nr_180_0 = 
        y_nr_enc[5] ^ 
        y_nr_enc[20] ^ 
        y_nr_enc[47] ^ 
0; ///1



    assign y_nr_p180 = 
y_nr_180_0 ^ 
0; ///3



wire y_nr_181_0;
assign y_nr_181_0 = 
        y_nr_enc[6] ^ 
        y_nr_enc[21] ^ 
        y_nr_enc[44] ^ 
0; ///1



    assign y_nr_p181 = 
y_nr_181_0 ^ 
0; ///3



wire y_nr_182_0;
assign y_nr_182_0 = 
        y_nr_enc[7] ^ 
        y_nr_enc[22] ^ 
        y_nr_enc[45] ^ 
0; ///1



    assign y_nr_p182 = 
y_nr_182_0 ^ 
0; ///3



wire y_nr_183_0;
assign y_nr_183_0 = 
        y_nr_enc[4] ^ 
        y_nr_enc[23] ^ 
        y_nr_enc[46] ^ 
0; ///1



    assign y_nr_p183 = 
y_nr_183_0 ^ 
0; ///3



wire y_nr_184_0;
assign y_nr_184_0 = 
        y_nr_enc[0] ^ 
        y_nr_enc[10] ^ 
        y_nr_enc[30] ^ 
0; ///1



    assign y_nr_p184 = 
y_nr_184_0 ^ 
0; ///3



wire y_nr_185_0;
assign y_nr_185_0 = 
        y_nr_enc[1] ^ 
        y_nr_enc[11] ^ 
        y_nr_enc[31] ^ 
0; ///1



    assign y_nr_p185 = 
y_nr_185_0 ^ 
0; ///3



wire y_nr_186_0;
assign y_nr_186_0 = 
        y_nr_enc[2] ^ 
        y_nr_enc[8] ^ 
        y_nr_enc[28] ^ 
0; ///1



    assign y_nr_p186 = 
y_nr_186_0 ^ 
0; ///3



wire y_nr_187_0;
assign y_nr_187_0 = 
        y_nr_enc[3] ^ 
        y_nr_enc[9] ^ 
        y_nr_enc[29] ^ 
0; ///1



    assign y_nr_p187 = 
y_nr_187_0 ^ 
0; ///3



wire y_nr_188_0;
assign y_nr_188_0 = 
        y_nr_enc[43] ^ 
        y_nr_enc[55] ^ 
0; ///1



    assign y_nr_p188 = 
y_nr_188_0 ^ 
0; ///3



wire y_nr_189_0;
assign y_nr_189_0 = 
        y_nr_enc[40] ^ 
        y_nr_enc[52] ^ 
0; ///1



    assign y_nr_p189 = 
y_nr_189_0 ^ 
0; ///3



wire y_nr_190_0;
assign y_nr_190_0 = 
        y_nr_enc[41] ^ 
        y_nr_enc[53] ^ 
0; ///1



    assign y_nr_p190 = 
y_nr_190_0 ^ 
0; ///3



wire y_nr_191_0;
assign y_nr_191_0 = 
        y_nr_enc[42] ^ 
        y_nr_enc[54] ^ 
0; ///1



    assign y_nr_p191 = 
y_nr_191_0 ^ 
0; ///3



wire y_nr_192_0;
assign y_nr_192_0 = 
        y_nr_enc[7] ^ 
        y_nr_enc[22] ^ 
        y_nr_enc[46] ^ 
0; ///1



    assign y_nr_p192 = 
y_nr_192_0 ^ 
0; ///3



wire y_nr_193_0;
assign y_nr_193_0 = 
        y_nr_enc[4] ^ 
        y_nr_enc[23] ^ 
        y_nr_enc[47] ^ 
0; ///1



    assign y_nr_p193 = 
y_nr_193_0 ^ 
0; ///3



wire y_nr_194_0;
assign y_nr_194_0 = 
        y_nr_enc[5] ^ 
        y_nr_enc[20] ^ 
        y_nr_enc[44] ^ 
0; ///1



    assign y_nr_p194 = 
y_nr_194_0 ^ 
0; ///3



wire y_nr_195_0;
assign y_nr_195_0 = 
        y_nr_enc[6] ^ 
        y_nr_enc[21] ^ 
        y_nr_enc[45] ^ 
0; ///1



    assign y_nr_p195 = 
y_nr_195_0 ^ 
0; ///3



wire y_nr_196_0;
assign y_nr_196_0 = 
        y_nr_enc[3] ^ 
        y_nr_enc[28] ^ 
        y_nr_enc[50] ^ 
0; ///1



    assign y_nr_p196 = 
y_nr_196_0 ^ 
0; ///3



wire y_nr_197_0;
assign y_nr_197_0 = 
        y_nr_enc[0] ^ 
        y_nr_enc[29] ^ 
        y_nr_enc[51] ^ 
0; ///1



    assign y_nr_p197 = 
y_nr_197_0 ^ 
0; ///3



wire y_nr_198_0;
assign y_nr_198_0 = 
        y_nr_enc[1] ^ 
        y_nr_enc[30] ^ 
        y_nr_enc[48] ^ 
0; ///1



    assign y_nr_p198 = 
y_nr_198_0 ^ 
0; ///3



wire y_nr_199_0;
assign y_nr_199_0 = 
        y_nr_enc[2] ^ 
        y_nr_enc[31] ^ 
        y_nr_enc[49] ^ 
0; ///1



    assign y_nr_p199 = 
y_nr_199_0 ^ 
0; ///3



wire y_nr_200_0;
assign y_nr_200_0 = 
        y_nr_enc[8] ^ 
        y_nr_enc[43] ^ 
        y_nr_enc[52] ^ 
0; ///1



    assign y_nr_p200 = 
y_nr_200_0 ^ 
0; ///3



wire y_nr_201_0;
assign y_nr_201_0 = 
        y_nr_enc[9] ^ 
        y_nr_enc[40] ^ 
        y_nr_enc[53] ^ 
0; ///1



    assign y_nr_p201 = 
y_nr_201_0 ^ 
0; ///3



wire y_nr_202_0;
assign y_nr_202_0 = 
        y_nr_enc[10] ^ 
        y_nr_enc[41] ^ 
        y_nr_enc[54] ^ 
0; ///1



    assign y_nr_p202 = 
y_nr_202_0 ^ 
0; ///3



wire y_nr_203_0;
assign y_nr_203_0 = 
        y_nr_enc[11] ^ 
        y_nr_enc[42] ^ 
        y_nr_enc[55] ^ 
0; ///1



    assign y_nr_p203 = 
y_nr_203_0 ^ 
0; ///3



wire y_nr_204_0;
assign y_nr_204_0 = 
        y_nr_enc[5] ^ 
        y_nr_enc[21] ^ 
        y_nr_enc[46] ^ 
0; ///1



    assign y_nr_p204 = 
y_nr_204_0 ^ 
0; ///3



wire y_nr_205_0;
assign y_nr_205_0 = 
        y_nr_enc[6] ^ 
        y_nr_enc[22] ^ 
        y_nr_enc[47] ^ 
0; ///1



    assign y_nr_p205 = 
y_nr_205_0 ^ 
0; ///3



wire y_nr_206_0;
assign y_nr_206_0 = 
        y_nr_enc[7] ^ 
        y_nr_enc[23] ^ 
        y_nr_enc[44] ^ 
0; ///1



    assign y_nr_p206 = 
y_nr_206_0 ^ 
0; ///3



wire y_nr_207_0;
assign y_nr_207_0 = 
        y_nr_enc[4] ^ 
        y_nr_enc[20] ^ 
        y_nr_enc[45] ^ 
0; ///1



    assign y_nr_p207 = 
y_nr_207_0 ^ 
0; ///3



