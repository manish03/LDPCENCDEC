reg [fgallag_WDTH -1:0] fgallag0x00002_0, fgallag0x00002_0_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_1, fgallag0x00002_1_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_2, fgallag0x00002_2_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_3, fgallag0x00002_3_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_4, fgallag0x00002_4_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_5, fgallag0x00002_5_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_6, fgallag0x00002_6_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_7, fgallag0x00002_7_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_8, fgallag0x00002_8_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_9, fgallag0x00002_9_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_10, fgallag0x00002_10_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_11, fgallag0x00002_11_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_12, fgallag0x00002_12_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_13, fgallag0x00002_13_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_14, fgallag0x00002_14_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_15, fgallag0x00002_15_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_16, fgallag0x00002_16_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_17, fgallag0x00002_17_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_18, fgallag0x00002_18_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_19, fgallag0x00002_19_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_20, fgallag0x00002_20_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_21, fgallag0x00002_21_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_22, fgallag0x00002_22_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_23, fgallag0x00002_23_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_24, fgallag0x00002_24_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_25, fgallag0x00002_25_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_26, fgallag0x00002_26_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_27, fgallag0x00002_27_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_28, fgallag0x00002_28_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_29, fgallag0x00002_29_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_30, fgallag0x00002_30_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_31, fgallag0x00002_31_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_32, fgallag0x00002_32_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_33, fgallag0x00002_33_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_34, fgallag0x00002_34_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_35, fgallag0x00002_35_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_36, fgallag0x00002_36_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_37, fgallag0x00002_37_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_38, fgallag0x00002_38_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_39, fgallag0x00002_39_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_40, fgallag0x00002_40_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_41, fgallag0x00002_41_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_42, fgallag0x00002_42_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_43, fgallag0x00002_43_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_44, fgallag0x00002_44_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_45, fgallag0x00002_45_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_46, fgallag0x00002_46_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_47, fgallag0x00002_47_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_48, fgallag0x00002_48_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_49, fgallag0x00002_49_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_50, fgallag0x00002_50_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_51, fgallag0x00002_51_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_52, fgallag0x00002_52_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_53, fgallag0x00002_53_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_54, fgallag0x00002_54_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_55, fgallag0x00002_55_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_56, fgallag0x00002_56_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_57, fgallag0x00002_57_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_58, fgallag0x00002_58_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_59, fgallag0x00002_59_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_60, fgallag0x00002_60_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_61, fgallag0x00002_61_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_62, fgallag0x00002_62_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_63, fgallag0x00002_63_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_64, fgallag0x00002_64_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_65, fgallag0x00002_65_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_66, fgallag0x00002_66_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_67, fgallag0x00002_67_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_68, fgallag0x00002_68_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_69, fgallag0x00002_69_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_70, fgallag0x00002_70_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_71, fgallag0x00002_71_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_72, fgallag0x00002_72_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_73, fgallag0x00002_73_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_74, fgallag0x00002_74_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_75, fgallag0x00002_75_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_76, fgallag0x00002_76_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_77, fgallag0x00002_77_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_78, fgallag0x00002_78_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_79, fgallag0x00002_79_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_80, fgallag0x00002_80_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_81, fgallag0x00002_81_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_82, fgallag0x00002_82_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_83, fgallag0x00002_83_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_84, fgallag0x00002_84_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_85, fgallag0x00002_85_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_86, fgallag0x00002_86_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_87, fgallag0x00002_87_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_88, fgallag0x00002_88_q;
reg [fgallag_WDTH -1:0] fgallag0x00002_89, fgallag0x00002_89_q;
reg start_d_fgallag0x00002_q ;
always_comb begin
 fgallag0x00002_0_q =  fgallag0x00002_0;
 fgallag0x00002_1_q =  fgallag0x00002_1;
 fgallag0x00002_2_q =  fgallag0x00002_2;
 fgallag0x00002_3_q =  fgallag0x00002_3;
 fgallag0x00002_4_q =  fgallag0x00002_4;
 fgallag0x00002_5_q =  fgallag0x00002_5;
 fgallag0x00002_6_q =  fgallag0x00002_6;
 fgallag0x00002_7_q =  fgallag0x00002_7;
 fgallag0x00002_8_q =  fgallag0x00002_8;
 fgallag0x00002_9_q =  fgallag0x00002_9;
 fgallag0x00002_10_q =  fgallag0x00002_10;
 fgallag0x00002_11_q =  fgallag0x00002_11;
 fgallag0x00002_12_q =  fgallag0x00002_12;
 fgallag0x00002_13_q =  fgallag0x00002_13;
 fgallag0x00002_14_q =  fgallag0x00002_14;
 fgallag0x00002_15_q =  fgallag0x00002_15;
 fgallag0x00002_16_q =  fgallag0x00002_16;
 fgallag0x00002_17_q =  fgallag0x00002_17;
 fgallag0x00002_18_q =  fgallag0x00002_18;
 fgallag0x00002_19_q =  fgallag0x00002_19;
 fgallag0x00002_20_q =  fgallag0x00002_20;
 fgallag0x00002_21_q =  fgallag0x00002_21;
 fgallag0x00002_22_q =  fgallag0x00002_22;
 fgallag0x00002_23_q =  fgallag0x00002_23;
 fgallag0x00002_24_q =  fgallag0x00002_24;
 fgallag0x00002_25_q =  fgallag0x00002_25;
 fgallag0x00002_26_q =  fgallag0x00002_26;
 fgallag0x00002_27_q =  fgallag0x00002_27;
 fgallag0x00002_28_q =  fgallag0x00002_28;
 fgallag0x00002_29_q =  fgallag0x00002_29;
 fgallag0x00002_30_q =  fgallag0x00002_30;
 fgallag0x00002_31_q =  fgallag0x00002_31;
 fgallag0x00002_32_q =  fgallag0x00002_32;
 fgallag0x00002_33_q =  fgallag0x00002_33;
 fgallag0x00002_34_q =  fgallag0x00002_34;
 fgallag0x00002_35_q =  fgallag0x00002_35;
 fgallag0x00002_36_q =  fgallag0x00002_36;
 fgallag0x00002_37_q =  fgallag0x00002_37;
 fgallag0x00002_38_q =  fgallag0x00002_38;
 fgallag0x00002_39_q =  fgallag0x00002_39;
 fgallag0x00002_40_q =  fgallag0x00002_40;
 fgallag0x00002_41_q =  fgallag0x00002_41;
 fgallag0x00002_42_q =  fgallag0x00002_42;
 fgallag0x00002_43_q =  fgallag0x00002_43;
 fgallag0x00002_44_q =  fgallag0x00002_44;
 fgallag0x00002_45_q =  fgallag0x00002_45;
 fgallag0x00002_46_q =  fgallag0x00002_46;
 fgallag0x00002_47_q =  fgallag0x00002_47;
 fgallag0x00002_48_q =  fgallag0x00002_48;
 fgallag0x00002_49_q =  fgallag0x00002_49;
 fgallag0x00002_50_q =  fgallag0x00002_50;
 fgallag0x00002_51_q =  fgallag0x00002_51;
 fgallag0x00002_52_q =  fgallag0x00002_52;
 fgallag0x00002_53_q =  fgallag0x00002_53;
 fgallag0x00002_54_q =  fgallag0x00002_54;
 fgallag0x00002_55_q =  fgallag0x00002_55;
 fgallag0x00002_56_q =  fgallag0x00002_56;
 fgallag0x00002_57_q =  fgallag0x00002_57;
 fgallag0x00002_58_q =  fgallag0x00002_58;
 fgallag0x00002_59_q =  fgallag0x00002_59;
 fgallag0x00002_60_q =  fgallag0x00002_60;
 fgallag0x00002_61_q =  fgallag0x00002_61;
 fgallag0x00002_62_q =  fgallag0x00002_62;
 fgallag0x00002_63_q =  fgallag0x00002_63;
 fgallag0x00002_64_q =  fgallag0x00002_64;
 fgallag0x00002_65_q =  fgallag0x00002_65;
 fgallag0x00002_66_q =  fgallag0x00002_66;
 fgallag0x00002_67_q =  fgallag0x00002_67;
 fgallag0x00002_68_q =  fgallag0x00002_68;
 fgallag0x00002_69_q =  fgallag0x00002_69;
 fgallag0x00002_70_q =  fgallag0x00002_70;
 fgallag0x00002_71_q =  fgallag0x00002_71;
 fgallag0x00002_72_q =  fgallag0x00002_72;
 fgallag0x00002_73_q =  fgallag0x00002_73;
 fgallag0x00002_74_q =  fgallag0x00002_74;
 fgallag0x00002_75_q =  fgallag0x00002_75;
 fgallag0x00002_76_q =  fgallag0x00002_76;
 fgallag0x00002_77_q =  fgallag0x00002_77;
 fgallag0x00002_78_q =  fgallag0x00002_78;
 fgallag0x00002_79_q =  fgallag0x00002_79;
 fgallag0x00002_80_q =  fgallag0x00002_80;
 fgallag0x00002_81_q =  fgallag0x00002_81;
 fgallag0x00002_82_q =  fgallag0x00002_82;
 fgallag0x00002_83_q =  fgallag0x00002_83;
 fgallag0x00002_84_q =  fgallag0x00002_84;
 fgallag0x00002_85_q =  fgallag0x00002_85;
 fgallag0x00002_86_q =  fgallag0x00002_86;
 fgallag0x00002_87_q =  fgallag0x00002_87;
 fgallag0x00002_88_q =  fgallag0x00002_88;
 fgallag0x00002_89_q =  fgallag0x00002_89;
 start_d_fgallag0x00002_q =  start_d_fgallag0x00001_q;
end
