              fgallag0x00004_0 = 
          (!fgallag_sel[3]) ? 
                       fgallag0x00003_0_q: 
                       fgallag0x00003_1_q;
              fgallag0x00004_1 = 
          (!fgallag_sel[3]) ? 
                       fgallag0x00003_2_q: 
                       fgallag0x00003_3_q;
              fgallag0x00004_2 = 
          (!fgallag_sel[3]) ? 
                       fgallag0x00003_4_q: 
                       fgallag0x00003_5_q;
              fgallag0x00004_3 = 
          (!fgallag_sel[3]) ? 
                       fgallag0x00003_6_q: 
                       fgallag0x00003_7_q;
              fgallag0x00004_4 = 
          (!fgallag_sel[3]) ? 
                       fgallag0x00003_8_q: 
                       fgallag0x00003_9_q;
              fgallag0x00004_5 = 
          (!fgallag_sel[3]) ? 
                       fgallag0x00003_10_q: 
                       fgallag0x00003_11_q;
              fgallag0x00004_6 = 
          (!fgallag_sel[3]) ? 
                       fgallag0x00003_12_q: 
                       fgallag0x00003_13_q;
              fgallag0x00004_7 = 
          (!fgallag_sel[3]) ? 
                       fgallag0x00003_14_q: 
                       fgallag0x00003_15_q;
              fgallag0x00004_8 = 
          (!fgallag_sel[3]) ? 
                       fgallag0x00003_16_q: 
                       fgallag0x00003_17_q;
              fgallag0x00004_9 = 
          (!fgallag_sel[3]) ? 
                       fgallag0x00003_18_q: 
                       fgallag0x00003_19_q;
              fgallag0x00004_10 = 
          (!fgallag_sel[3]) ? 
                       fgallag0x00003_20_q: 
                       fgallag0x00003_21_q;
              fgallag0x00004_11 = 
          (!fgallag_sel[3]) ? 
                       fgallag0x00003_22_q: 
                       fgallag0x00003_23_q;
              fgallag0x00004_12 = 
          (!fgallag_sel[3]) ? 
                       fgallag0x00003_24_q: 
                       fgallag0x00003_25_q;
              fgallag0x00004_13 = 
          (!fgallag_sel[3]) ? 
                       fgallag0x00003_26_q: 
                       fgallag0x00003_27_q;
              fgallag0x00004_14 = 
          (!fgallag_sel[3]) ? 
                       fgallag0x00003_28_q: 
                       fgallag0x00003_29_q;
              fgallag0x00004_15 = 
          (!fgallag_sel[3]) ? 
                       fgallag0x00003_30_q: 
                       fgallag0x00003_31_q;
               fgallag0x00004_16 =  fgallag0x00003_32_q ;
              fgallag0x00004_17 = 
          (!fgallag_sel[3]) ? 
                       fgallag0x00003_34_q: 
                       fgallag0x00003_35_q;
               fgallag0x00004_18 =  fgallag0x00003_36_q ;
               fgallag0x00004_19 =  fgallag0x00003_38_q ;
               fgallag0x00004_20 =  fgallag0x00003_40_q ;
               fgallag0x00004_21 =  fgallag0x00003_42_q ;
              fgallag0x00004_22 = 
          (!fgallag_sel[3]) ? 
                       fgallag0x00003_44_q: 
                       fgallag0x00003_45_q;
               fgallag0x00004_23 =  0;
