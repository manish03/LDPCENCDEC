              flogtanh0x00003_0 = 
          (!flogtanh_sel[2]) ? 
                       flogtanh0x00002_0_q: 
                       flogtanh0x00002_1_q;
              flogtanh0x00003_1 = 
          (!flogtanh_sel[2]) ? 
                       flogtanh0x00002_2_q: 
                       flogtanh0x00002_3_q;
              flogtanh0x00003_2 = 
          (!flogtanh_sel[2]) ? 
                       flogtanh0x00002_4_q: 
                       flogtanh0x00002_5_q;
              flogtanh0x00003_3 = 
          (!flogtanh_sel[2]) ? 
                       flogtanh0x00002_6_q: 
                       flogtanh0x00002_7_q;
              flogtanh0x00003_4 = 
          (!flogtanh_sel[2]) ? 
                       flogtanh0x00002_8_q: 
                       flogtanh0x00002_9_q;
              flogtanh0x00003_5 = 
          (!flogtanh_sel[2]) ? 
                       flogtanh0x00002_10_q: 
                       flogtanh0x00002_11_q;
              flogtanh0x00003_6 = 
          (!flogtanh_sel[2]) ? 
                       flogtanh0x00002_12_q: 
                       flogtanh0x00002_13_q;
              flogtanh0x00003_7 = 
          (!flogtanh_sel[2]) ? 
                       flogtanh0x00002_14_q: 
                       flogtanh0x00002_15_q;
              flogtanh0x00003_8 = 
          (!flogtanh_sel[2]) ? 
                       flogtanh0x00002_16_q: 
                       flogtanh0x00002_17_q;
              flogtanh0x00003_9 = 
          (!flogtanh_sel[2]) ? 
                       flogtanh0x00002_18_q: 
                       flogtanh0x00002_19_q;
              flogtanh0x00003_10 = 
          (!flogtanh_sel[2]) ? 
                       flogtanh0x00002_20_q: 
                       flogtanh0x00002_21_q;
              flogtanh0x00003_11 = 
          (!flogtanh_sel[2]) ? 
                       flogtanh0x00002_22_q: 
                       flogtanh0x00002_23_q;
              flogtanh0x00003_12 = 
          (!flogtanh_sel[2]) ? 
                       flogtanh0x00002_24_q: 
                       flogtanh0x00002_25_q;
              flogtanh0x00003_13 = 
          (!flogtanh_sel[2]) ? 
                       flogtanh0x00002_26_q: 
                       flogtanh0x00002_27_q;
              flogtanh0x00003_14 = 
          (!flogtanh_sel[2]) ? 
                       flogtanh0x00002_28_q: 
                       flogtanh0x00002_29_q;
              flogtanh0x00003_15 = 
          (!flogtanh_sel[2]) ? 
                       flogtanh0x00002_30_q: 
                       flogtanh0x00002_31_q;
              flogtanh0x00003_16 = 
          (!flogtanh_sel[2]) ? 
                       flogtanh0x00002_32_q: 
                       flogtanh0x00002_33_q;
              flogtanh0x00003_17 = 
          (!flogtanh_sel[2]) ? 
                       flogtanh0x00002_34_q: 
                       flogtanh0x00002_35_q;
              flogtanh0x00003_18 = 
          (!flogtanh_sel[2]) ? 
                       flogtanh0x00002_36_q: 
                       flogtanh0x00002_37_q;
              flogtanh0x00003_19 = 
          (!flogtanh_sel[2]) ? 
                       flogtanh0x00002_38_q: 
                       flogtanh0x00002_39_q;
              flogtanh0x00003_20 = 
          (!flogtanh_sel[2]) ? 
                       flogtanh0x00002_40_q: 
                       flogtanh0x00002_41_q;
              flogtanh0x00003_21 = 
          (!flogtanh_sel[2]) ? 
                       flogtanh0x00002_42_q: 
                       flogtanh0x00002_43_q;
              flogtanh0x00003_22 = 
          (!flogtanh_sel[2]) ? 
                       flogtanh0x00002_44_q: 
                       flogtanh0x00002_45_q;
              flogtanh0x00003_23 = 
          (!flogtanh_sel[2]) ? 
                       flogtanh0x00002_46_q: 
                       flogtanh0x00002_47_q;
               flogtanh0x00003_24 =  flogtanh0x00002_48_q ;
              flogtanh0x00003_25 = 
          (!flogtanh_sel[2]) ? 
                       flogtanh0x00002_50_q: 
                       flogtanh0x00002_51_q;
              flogtanh0x00003_26 = 
          (!flogtanh_sel[2]) ? 
                       flogtanh0x00002_52_q: 
                       flogtanh0x00002_53_q;
               flogtanh0x00003_27 =  flogtanh0x00002_54_q ;
              flogtanh0x00003_28 = 
          (!flogtanh_sel[2]) ? 
                       flogtanh0x00002_56_q: 
                       flogtanh0x00002_57_q;
               flogtanh0x00003_29 =  flogtanh0x00002_58_q ;
               flogtanh0x00003_30 =  flogtanh0x00002_60_q ;
              flogtanh0x00003_31 = 
          (!flogtanh_sel[2]) ? 
                       flogtanh0x00002_62_q: 
                       flogtanh0x00002_63_q;
               flogtanh0x00003_32 =  flogtanh0x00002_64_q ;
               flogtanh0x00003_33 =  flogtanh0x00002_66_q ;
               flogtanh0x00003_34 =  flogtanh0x00002_68_q ;
              flogtanh0x00003_35 = 
          (!flogtanh_sel[2]) ? 
                       flogtanh0x00002_70_q: 
                       flogtanh0x00002_71_q;
               flogtanh0x00003_36 =  flogtanh0x00002_72_q ;
               flogtanh0x00003_37 =  flogtanh0x00002_74_q ;
               flogtanh0x00003_38 =  flogtanh0x00002_76_q ;
               flogtanh0x00003_39 =  flogtanh0x00002_78_q ;
               flogtanh0x00003_40 =  flogtanh0x00002_80_q ;
               flogtanh0x00003_41 =  flogtanh0x00002_82_q ;
               flogtanh0x00003_42 =  flogtanh0x00002_84_q ;
               flogtanh0x00003_43 =  flogtanh0x00002_86_q ;
              flogtanh0x00003_44 = 
          (!flogtanh_sel[2]) ? 
                       flogtanh0x00002_88_q: 
                       flogtanh0x00002_89_q;
               flogtanh0x00003_45 =  0;
