              fgallag0xffffffff_0 = 
          (!fgallag_sel[8]) ? 
                       fgallag0x00008_0_q: 
                       fgallag0x00008_1_q;
               fgallag0xffffffff_1 =  0;
