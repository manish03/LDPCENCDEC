         fgallag0x00000_0 =   'h00380 ;
         fgallag0x00000_1 =   'h0013a ;
         fgallag0x00000_2 =   'h0011c ;
         fgallag0x00000_3 =   'h000fa ;
         fgallag0x00000_4 =   'h000e4 ;
         fgallag0x00000_5 =   'h000d4 ;
         fgallag0x00000_6 =   'h000c8 ;
         fgallag0x00000_7 =   'h000bd ;
         fgallag0x00000_8 =   'h000b4 ;
         fgallag0x00000_9 =   'h000ad ;
         fgallag0x00000_10 =   'h000a6 ;
         fgallag0x00000_11 =   'h0009f ;
         fgallag0x00000_12 =   'h0009a ;
         fgallag0x00000_13 =   'h00094 ;
         fgallag0x00000_14 =   'h0008f ;
         fgallag0x00000_15 =   'h0008b ;
         fgallag0x00000_16 =   'h00087 ;
         fgallag0x00000_17 =   'h00083 ;
         fgallag0x00000_18 =   'h0007f ;
         fgallag0x00000_19 =   'h0007c ;
         fgallag0x00000_20 =   'h00078 ;
         fgallag0x00000_21 =   'h00075 ;
         fgallag0x00000_22 =   'h00072 ;
         fgallag0x00000_23 =   'h0006f ;
         fgallag0x00000_24 =   'h0006d ;
         fgallag0x00000_25 =   'h0006a ;
         fgallag0x00000_26 =   'h00068 ;
         fgallag0x00000_27 =   'h00065 ;
         fgallag0x00000_28 =   'h00063 ;
         fgallag0x00000_29 =   'h00061 ;
         fgallag0x00000_30 =   'h0005f ;
         fgallag0x00000_31 =   'h0005d ;
         fgallag0x00000_32 =   'h0005b ;
         fgallag0x00000_33 =   'h00059 ;
         fgallag0x00000_34 =   'h00057 ;
         fgallag0x00000_35 =   'h00055 ;
         fgallag0x00000_36 =   'h00053 ;
         fgallag0x00000_37 =   'h00052 ;
         fgallag0x00000_38 =   'h00050 ;
         fgallag0x00000_39 =   'h0004f ;
         fgallag0x00000_40 =   'h0004d ;
         fgallag0x00000_41 =   'h0004b ;
         fgallag0x00000_42 =   'h0004a ;
         fgallag0x00000_43 =   'h00049 ;
         fgallag0x00000_44 =   'h00047 ;
         fgallag0x00000_45 =   'h00046 ;
         fgallag0x00000_46 =   'h00045 ;
         fgallag0x00000_47 =   'h00043 ;
         fgallag0x00000_48 =   'h00042 ;
         fgallag0x00000_49 =   'h00041 ;
         fgallag0x00000_50 =   'h00040 ;
         fgallag0x00000_51 =   'h0003f ;
         fgallag0x00000_52 =   'h0003d ;
         fgallag0x00000_53 =   'h0003c ;
         fgallag0x00000_54 =   'h0003b ;
         fgallag0x00000_55 =   'h0003a ;
         fgallag0x00000_56 =   'h00039 ;
         fgallag0x00000_57 =   'h00038 ;
         fgallag0x00000_58 =   'h00037 ;
         fgallag0x00000_59 =   'h00036 ;
         fgallag0x00000_60 =   'h00035 ;
         fgallag0x00000_61 =   'h00034 ;
         fgallag0x00000_62 =   'h00033 ;
         fgallag0x00000_63 =   'h00033 ;
         fgallag0x00000_64 =   'h00032 ;
         fgallag0x00000_65 =   'h00031 ;
         fgallag0x00000_66 =   'h00030 ;
         fgallag0x00000_67 =   'h0002f ;
         fgallag0x00000_68 =   'h0002e ;
         fgallag0x00000_69 =   'h0002e ;
         fgallag0x00000_70 =   'h0002d ;
         fgallag0x00000_71 =   'h0002c ;
         fgallag0x00000_72 =   'h0002b ;
         fgallag0x00000_73 =   'h0002b ;
         fgallag0x00000_74 =   'h0002a ;
         fgallag0x00000_75 =   'h00029 ;
         fgallag0x00000_76 =   'h00029 ;
         fgallag0x00000_77 =   'h00028 ;
         fgallag0x00000_78 =   'h00027 ;
         fgallag0x00000_79 =   'h00027 ;
         fgallag0x00000_80 =   'h00026 ;
         fgallag0x00000_81 =   'h00025 ;
         fgallag0x00000_82 =   'h00025 ;
         fgallag0x00000_83 =   'h00024 ;
         fgallag0x00000_84 =   'h00024 ;
         fgallag0x00000_85 =   'h00023 ;
         fgallag0x00000_86 =   'h00022 ;
         fgallag0x00000_87 =   'h00022 ;
         fgallag0x00000_88 =   'h00021 ;
         fgallag0x00000_89 =   'h00021 ;
         fgallag0x00000_90 =   'h00020 ;
         fgallag0x00000_91 =   'h00020 ;
         fgallag0x00000_92 =   'h0001f ;
         fgallag0x00000_93 =   'h0001f ;
         fgallag0x00000_94 =   'h0001e ;
         fgallag0x00000_95 =   'h0001e ;
         fgallag0x00000_96 =   'h0001d ;
         fgallag0x00000_97 =   'h0001d ;
         fgallag0x00000_98 =   'h0001c ;
         fgallag0x00000_99 =   'h0001c ;
         fgallag0x00000_100 =   'h0001b ;
         fgallag0x00000_101 =   'h0001b ;
         fgallag0x00000_102 =   'h0001b ;
         fgallag0x00000_103 =   'h0001a ;
         fgallag0x00000_104 =   'h0001a ;
         fgallag0x00000_105 =   'h00019 ;
         fgallag0x00000_106 =   'h00019 ;
         fgallag0x00000_107 =   'h00018 ;
         fgallag0x00000_108 =   'h00018 ;
         fgallag0x00000_109 =   'h00018 ;
         fgallag0x00000_110 =   'h00017 ;
         fgallag0x00000_111 =   'h00017 ;
         fgallag0x00000_112 =   'h00017 ;
         fgallag0x00000_113 =   'h00016 ;
         fgallag0x00000_114 =   'h00016 ;
         fgallag0x00000_115 =   'h00016 ;
         fgallag0x00000_116 =   'h00015 ;
         fgallag0x00000_117 =   'h00015 ;
         fgallag0x00000_118 =   'h00015 ;
         fgallag0x00000_119 =   'h00014 ;
         fgallag0x00000_120 =   'h00014 ;
         fgallag0x00000_121 =   'h00014 ;
         fgallag0x00000_122 =   'h00013 ;
         fgallag0x00000_123 =   'h00013 ;
         fgallag0x00000_124 =   'h00013 ;
         fgallag0x00000_125 =   'h00012 ;
         fgallag0x00000_126 =   'h00012 ;
         fgallag0x00000_127 =   'h00012 ;
         fgallag0x00000_128 =   'h00012 ;
         fgallag0x00000_129 =   'h00011 ;
         fgallag0x00000_130 =   'h00011 ;
         fgallag0x00000_131 =   'h00011 ;
         fgallag0x00000_132 =   'h00010 ;
         fgallag0x00000_133 =   'h00010 ;
         fgallag0x00000_134 =   'h00010 ;
         fgallag0x00000_135 =   'h00010 ;
         fgallag0x00000_136 =   'h0000f ;
         fgallag0x00000_137 =   'h0000f ;
         fgallag0x00000_138 =   'h0000f ;
         fgallag0x00000_139 =   'h0000f ;
         fgallag0x00000_140 =   'h0000e ;
         fgallag0x00000_141 =   'h0000e ;
         fgallag0x00000_142 =   'h0000e ;
         fgallag0x00000_143 =   'h0000e ;
         fgallag0x00000_144 =   'h0000e ;
         fgallag0x00000_145 =   'h0000d ;
         fgallag0x00000_146 =   'h0000d ;
         fgallag0x00000_147 =   'h0000d ;
         fgallag0x00000_148 =   'h0000d ;
         fgallag0x00000_149 =   'h0000d ;
         fgallag0x00000_150 =   'h0000c ;
         fgallag0x00000_151 =   'h0000c ;
         fgallag0x00000_152 =   'h0000c ;
         fgallag0x00000_153 =   'h0000c ;
         fgallag0x00000_154 =   'h0000c ;
         fgallag0x00000_155 =   'h0000b ;
         fgallag0x00000_156 =   'h0000b ;
         fgallag0x00000_157 =   'h0000b ;
         fgallag0x00000_158 =   'h0000b ;
         fgallag0x00000_159 =   'h0000b ;
         fgallag0x00000_160 =   'h0000b ;
         fgallag0x00000_161 =   'h0000a ;
         fgallag0x00000_162 =   'h0000a ;
         fgallag0x00000_163 =   'h0000a ;
         fgallag0x00000_164 =   'h0000a ;
         fgallag0x00000_165 =   'h0000a ;
         fgallag0x00000_166 =   'h0000a ;
         fgallag0x00000_167 =   'h00009 ;
         fgallag0x00000_168 =   'h00009 ;
         fgallag0x00000_169 =   'h00009 ;
         fgallag0x00000_170 =   'h00009 ;
         fgallag0x00000_171 =   'h00009 ;
         fgallag0x00000_172 =   'h00009 ;
         fgallag0x00000_173 =   'h00009 ;
         fgallag0x00000_174 =   'h00008 ;
         fgallag0x00000_175 =   'h00008 ;
         fgallag0x00000_176 =   'h00008 ;
         fgallag0x00000_177 =   'h00008 ;
         fgallag0x00000_178 =   'h00008 ;
         fgallag0x00000_179 =   'h00008 ;
         fgallag0x00000_180 =   'h00008 ;
         fgallag0x00000_181 =   'h00008 ;
         fgallag0x00000_182 =   'h00007 ;
         fgallag0x00000_183 =   'h00007 ;
         fgallag0x00000_184 =   'h00007 ;
         fgallag0x00000_185 =   'h00007 ;
         fgallag0x00000_186 =   'h00007 ;
         fgallag0x00000_187 =   'h00007 ;
         fgallag0x00000_188 =   'h00007 ;
         fgallag0x00000_189 =   'h00007 ;
         fgallag0x00000_190 =   'h00007 ;
         fgallag0x00000_191 =   'h00007 ;
         fgallag0x00000_192 =   'h00006 ;
         fgallag0x00000_193 =   'h00006 ;
         fgallag0x00000_194 =   'h00006 ;
         fgallag0x00000_195 =   'h00006 ;
         fgallag0x00000_196 =   'h00006 ;
         fgallag0x00000_197 =   'h00006 ;
         fgallag0x00000_198 =   'h00006 ;
         fgallag0x00000_199 =   'h00006 ;
         fgallag0x00000_200 =   'h00006 ;
         fgallag0x00000_201 =   'h00006 ;
         fgallag0x00000_202 =   'h00005 ;
         fgallag0x00000_203 =   'h00005 ;
         fgallag0x00000_204 =   'h00005 ;
         fgallag0x00000_205 =   'h00005 ;
         fgallag0x00000_206 =   'h00005 ;
         fgallag0x00000_207 =   'h00005 ;
         fgallag0x00000_208 =   'h00005 ;
         fgallag0x00000_209 =   'h00005 ;
         fgallag0x00000_210 =   'h00005 ;
         fgallag0x00000_211 =   'h00005 ;
         fgallag0x00000_212 =   'h00005 ;
         fgallag0x00000_213 =   'h00005 ;
         fgallag0x00000_214 =   'h00005 ;
         fgallag0x00000_215 =   'h00004 ;
         fgallag0x00000_216 =   'h00004 ;
         fgallag0x00000_217 =   'h00004 ;
         fgallag0x00000_218 =   'h00004 ;
         fgallag0x00000_219 =   'h00004 ;
         fgallag0x00000_220 =   'h00004 ;
         fgallag0x00000_221 =   'h00004 ;
         fgallag0x00000_222 =   'h00004 ;
         fgallag0x00000_223 =   'h00004 ;
         fgallag0x00000_224 =   'h00004 ;
         fgallag0x00000_225 =   'h00004 ;
         fgallag0x00000_226 =   'h00004 ;
         fgallag0x00000_227 =   'h00004 ;
         fgallag0x00000_228 =   'h00004 ;
         fgallag0x00000_229 =   'h00004 ;
         fgallag0x00000_230 =   'h00004 ;
         fgallag0x00000_231 =   'h00003 ;
         fgallag0x00000_232 =   'h00003 ;
         fgallag0x00000_233 =   'h00003 ;
         fgallag0x00000_234 =   'h00003 ;
         fgallag0x00000_235 =   'h00003 ;
         fgallag0x00000_236 =   'h00003 ;
         fgallag0x00000_237 =   'h00003 ;
         fgallag0x00000_238 =   'h00003 ;
         fgallag0x00000_239 =   'h00003 ;
         fgallag0x00000_240 =   'h00003 ;
         fgallag0x00000_241 =   'h00003 ;
         fgallag0x00000_242 =   'h00003 ;
         fgallag0x00000_243 =   'h00003 ;
         fgallag0x00000_244 =   'h00003 ;
         fgallag0x00000_245 =   'h00003 ;
         fgallag0x00000_246 =   'h00003 ;
         fgallag0x00000_247 =   'h00003 ;
         fgallag0x00000_248 =   'h00003 ;
         fgallag0x00000_249 =   'h00003 ;
         fgallag0x00000_250 =   'h00003 ;
         fgallag0x00000_251 =   'h00003 ;
         fgallag0x00000_252 =   'h00003 ;
         fgallag0x00000_253 =   'h00002 ;
         fgallag0x00000_254 =   'h00002 ;
         fgallag0x00000_255 =   'h00002 ;
         fgallag0x00000_256 =   'h00002 ;
         fgallag0x00000_257 =   'h00002 ;
         fgallag0x00000_258 =   'h00002 ;
         fgallag0x00000_259 =   'h00002 ;
         fgallag0x00000_260 =   'h00002 ;
         fgallag0x00000_261 =   'h00002 ;
         fgallag0x00000_262 =   'h00002 ;
         fgallag0x00000_263 =   'h00002 ;
         fgallag0x00000_264 =   'h00002 ;
         fgallag0x00000_265 =   'h00002 ;
         fgallag0x00000_266 =   'h00002 ;
         fgallag0x00000_267 =   'h00002 ;
         fgallag0x00000_268 =   'h00002 ;
         fgallag0x00000_269 =   'h00002 ;
         fgallag0x00000_270 =   'h00002 ;
         fgallag0x00000_271 =   'h00002 ;
         fgallag0x00000_272 =   'h00002 ;
         fgallag0x00000_273 =   'h00002 ;
         fgallag0x00000_274 =   'h00002 ;
         fgallag0x00000_275 =   'h00002 ;
         fgallag0x00000_276 =   'h00002 ;
         fgallag0x00000_277 =   'h00002 ;
         fgallag0x00000_278 =   'h00002 ;
         fgallag0x00000_279 =   'h00002 ;
         fgallag0x00000_280 =   'h00002 ;
         fgallag0x00000_281 =   'h00002 ;
         fgallag0x00000_282 =   'h00002 ;
         fgallag0x00000_283 =   'h00002 ;
         fgallag0x00000_284 =   'h00002 ;
         fgallag0x00000_285 =   'h00001 ;
         fgallag0x00000_286 =   'h00001 ;
         fgallag0x00000_287 =   'h00001 ;
         fgallag0x00000_288 =   'h00001 ;
         fgallag0x00000_289 =   'h00001 ;
         fgallag0x00000_290 =   'h00001 ;
         fgallag0x00000_291 =   'h00001 ;
         fgallag0x00000_292 =   'h00001 ;
         fgallag0x00000_293 =   'h00001 ;
         fgallag0x00000_294 =   'h00001 ;
         fgallag0x00000_295 =   'h00001 ;
         fgallag0x00000_296 =   'h00001 ;
         fgallag0x00000_297 =   'h00001 ;
         fgallag0x00000_298 =   'h00001 ;
         fgallag0x00000_299 =   'h00001 ;
         fgallag0x00000_300 =   'h00001 ;
         fgallag0x00000_301 =   'h00001 ;
         fgallag0x00000_302 =   'h00001 ;
         fgallag0x00000_303 =   'h00001 ;
         fgallag0x00000_304 =   'h00001 ;
         fgallag0x00000_305 =   'h00001 ;
         fgallag0x00000_306 =   'h00001 ;
         fgallag0x00000_307 =   'h00001 ;
         fgallag0x00000_308 =   'h00001 ;
         fgallag0x00000_309 =   'h00001 ;
         fgallag0x00000_310 =   'h00001 ;
         fgallag0x00000_311 =   'h00001 ;
         fgallag0x00000_312 =   'h00001 ;
         fgallag0x00000_313 =   'h00001 ;
         fgallag0x00000_314 =   'h00001 ;
         fgallag0x00000_315 =   'h00001 ;
         fgallag0x00000_316 =   'h00001 ;
         fgallag0x00000_317 =   'h00001 ;
         fgallag0x00000_318 =   'h00001 ;
         fgallag0x00000_319 =   'h00001 ;
         fgallag0x00000_320 =   'h00001 ;
         fgallag0x00000_321 =   'h00001 ;
         fgallag0x00000_322 =   'h00001 ;
         fgallag0x00000_323 =   'h00001 ;
         fgallag0x00000_324 =   'h00001 ;
         fgallag0x00000_325 =   'h00001 ;
         fgallag0x00000_326 =   'h00001 ;
         fgallag0x00000_327 =   'h00001 ;
         fgallag0x00000_328 =   'h00001 ;
         fgallag0x00000_329 =   'h00001 ;
         fgallag0x00000_330 =   'h00001 ;
         fgallag0x00000_331 =   'h00001 ;
         fgallag0x00000_332 =   'h00001 ;
         fgallag0x00000_333 =   'h00001 ;
         fgallag0x00000_334 =   'h00001 ;
         fgallag0x00000_335 =   'h00001 ;
         fgallag0x00000_336 =   'h00001 ;
         fgallag0x00000_337 =   'h00001 ;
         fgallag0x00000_338 =   'h00001 ;
         fgallag0x00000_339 =   'h00001 ;
         fgallag0x00000_340 =   'h00001 ;
         fgallag0x00000_341 =   'h00001 ;
         fgallag0x00000_342 =   'h00001 ;
         fgallag0x00000_343 =   'h00001 ;
         fgallag0x00000_344 =   'h00001 ;
         fgallag0x00000_345 =   'h00001 ;
         fgallag0x00000_346 =   'h00001 ;
         fgallag0x00000_347 =   'h00001 ;
         fgallag0x00000_348 =   'h00001 ;
         fgallag0x00000_349 =   'h00001 ;
         fgallag0x00000_350 =   'h00001 ;
         fgallag0x00000_351 =   'h00001 ;
         fgallag0x00000_352 =   'h00001 ;
         fgallag0x00000_353 =   'h00001 ;
         fgallag0x00000_354 =   'h00001 ;
         fgallag0x00000_355 =   'h00001 ;
