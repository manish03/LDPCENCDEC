package LDPC_CSR_rtl_pkg;
  localparam int LDPC_ENC_MSG_IN_0_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_0_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_0_BYTE_OFFSET = 13'h0000;
  localparam int LDPC_ENC_MSG_IN_0_MSG_IN_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_0_MSG_IN_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_0_MSG_IN_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_1_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_1_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_1_BYTE_OFFSET = 13'h0004;
  localparam int LDPC_ENC_MSG_IN_1_MSG_IN_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_1_MSG_IN_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_1_MSG_IN_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_2_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_2_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_2_BYTE_OFFSET = 13'h0008;
  localparam int LDPC_ENC_MSG_IN_2_MSG_IN_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_2_MSG_IN_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_2_MSG_IN_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_3_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_3_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_3_BYTE_OFFSET = 13'h000c;
  localparam int LDPC_ENC_MSG_IN_3_MSG_IN_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_3_MSG_IN_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_3_MSG_IN_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_4_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_4_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_4_BYTE_OFFSET = 13'h0010;
  localparam int LDPC_ENC_MSG_IN_4_MSG_IN_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_4_MSG_IN_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_4_MSG_IN_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_5_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_5_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_5_BYTE_OFFSET = 13'h0014;
  localparam int LDPC_ENC_MSG_IN_5_MSG_IN_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_5_MSG_IN_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_5_MSG_IN_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_6_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_6_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_6_BYTE_OFFSET = 13'h0018;
  localparam int LDPC_ENC_MSG_IN_6_MSG_IN_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_6_MSG_IN_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_6_MSG_IN_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_7_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_7_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_7_BYTE_OFFSET = 13'h001c;
  localparam int LDPC_ENC_MSG_IN_7_MSG_IN_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_7_MSG_IN_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_7_MSG_IN_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_8_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_8_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_8_BYTE_OFFSET = 13'h0020;
  localparam int LDPC_ENC_MSG_IN_8_MSG_IN_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_8_MSG_IN_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_8_MSG_IN_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_9_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_9_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_9_BYTE_OFFSET = 13'h0024;
  localparam int LDPC_ENC_MSG_IN_9_MSG_IN_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_9_MSG_IN_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_9_MSG_IN_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_10_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_10_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_10_BYTE_OFFSET = 13'h0028;
  localparam int LDPC_ENC_MSG_IN_10_MSG_IN_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_10_MSG_IN_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_10_MSG_IN_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_11_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_11_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_11_BYTE_OFFSET = 13'h002c;
  localparam int LDPC_ENC_MSG_IN_11_MSG_IN_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_11_MSG_IN_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_11_MSG_IN_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_12_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_12_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_12_BYTE_OFFSET = 13'h0030;
  localparam int LDPC_ENC_MSG_IN_12_MSG_IN_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_12_MSG_IN_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_12_MSG_IN_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_13_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_13_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_13_BYTE_OFFSET = 13'h0034;
  localparam int LDPC_ENC_MSG_IN_13_MSG_IN_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_13_MSG_IN_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_13_MSG_IN_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_14_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_14_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_14_BYTE_OFFSET = 13'h0038;
  localparam int LDPC_ENC_MSG_IN_14_MSG_IN_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_14_MSG_IN_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_14_MSG_IN_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_15_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_15_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_15_BYTE_OFFSET = 13'h003c;
  localparam int LDPC_ENC_MSG_IN_15_MSG_IN_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_15_MSG_IN_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_15_MSG_IN_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_16_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_16_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_16_BYTE_OFFSET = 13'h0040;
  localparam int LDPC_ENC_MSG_IN_16_MSG_IN_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_16_MSG_IN_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_16_MSG_IN_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_17_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_17_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_17_BYTE_OFFSET = 13'h0044;
  localparam int LDPC_ENC_MSG_IN_17_MSG_IN_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_17_MSG_IN_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_17_MSG_IN_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_18_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_18_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_18_BYTE_OFFSET = 13'h0048;
  localparam int LDPC_ENC_MSG_IN_18_MSG_IN_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_18_MSG_IN_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_18_MSG_IN_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_19_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_19_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_19_BYTE_OFFSET = 13'h004c;
  localparam int LDPC_ENC_MSG_IN_19_MSG_IN_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_19_MSG_IN_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_19_MSG_IN_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_20_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_20_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_20_BYTE_OFFSET = 13'h0050;
  localparam int LDPC_ENC_MSG_IN_20_MSG_IN_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_20_MSG_IN_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_20_MSG_IN_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_21_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_21_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_21_BYTE_OFFSET = 13'h0054;
  localparam int LDPC_ENC_MSG_IN_21_MSG_IN_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_21_MSG_IN_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_21_MSG_IN_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_22_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_22_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_22_BYTE_OFFSET = 13'h0058;
  localparam int LDPC_ENC_MSG_IN_22_MSG_IN_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_22_MSG_IN_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_22_MSG_IN_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_23_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_23_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_23_BYTE_OFFSET = 13'h005c;
  localparam int LDPC_ENC_MSG_IN_23_MSG_IN_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_23_MSG_IN_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_23_MSG_IN_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_24_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_24_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_24_BYTE_OFFSET = 13'h0060;
  localparam int LDPC_ENC_MSG_IN_24_MSG_IN_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_24_MSG_IN_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_24_MSG_IN_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_25_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_25_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_25_BYTE_OFFSET = 13'h0064;
  localparam int LDPC_ENC_MSG_IN_25_MSG_IN_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_25_MSG_IN_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_25_MSG_IN_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_26_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_26_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_26_BYTE_OFFSET = 13'h0068;
  localparam int LDPC_ENC_MSG_IN_26_MSG_IN_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_26_MSG_IN_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_26_MSG_IN_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_27_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_27_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_27_BYTE_OFFSET = 13'h006c;
  localparam int LDPC_ENC_MSG_IN_27_MSG_IN_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_27_MSG_IN_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_27_MSG_IN_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_28_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_28_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_28_BYTE_OFFSET = 13'h0070;
  localparam int LDPC_ENC_MSG_IN_28_MSG_IN_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_28_MSG_IN_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_28_MSG_IN_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_29_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_29_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_29_BYTE_OFFSET = 13'h0074;
  localparam int LDPC_ENC_MSG_IN_29_MSG_IN_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_29_MSG_IN_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_29_MSG_IN_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_30_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_30_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_30_BYTE_OFFSET = 13'h0078;
  localparam int LDPC_ENC_MSG_IN_30_MSG_IN_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_30_MSG_IN_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_30_MSG_IN_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_31_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_31_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_31_BYTE_OFFSET = 13'h007c;
  localparam int LDPC_ENC_MSG_IN_31_MSG_IN_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_31_MSG_IN_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_31_MSG_IN_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_32_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_32_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_32_BYTE_OFFSET = 13'h0080;
  localparam int LDPC_ENC_MSG_IN_32_MSG_IN_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_32_MSG_IN_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_32_MSG_IN_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_33_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_33_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_33_BYTE_OFFSET = 13'h0084;
  localparam int LDPC_ENC_MSG_IN_33_MSG_IN_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_33_MSG_IN_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_33_MSG_IN_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_34_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_34_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_34_BYTE_OFFSET = 13'h0088;
  localparam int LDPC_ENC_MSG_IN_34_MSG_IN_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_34_MSG_IN_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_34_MSG_IN_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_35_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_35_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_35_BYTE_OFFSET = 13'h008c;
  localparam int LDPC_ENC_MSG_IN_35_MSG_IN_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_35_MSG_IN_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_35_MSG_IN_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_36_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_36_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_36_BYTE_OFFSET = 13'h0090;
  localparam int LDPC_ENC_MSG_IN_36_MSG_IN_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_36_MSG_IN_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_36_MSG_IN_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_37_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_37_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_37_BYTE_OFFSET = 13'h0094;
  localparam int LDPC_ENC_MSG_IN_37_MSG_IN_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_37_MSG_IN_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_37_MSG_IN_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_38_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_38_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_38_BYTE_OFFSET = 13'h0098;
  localparam int LDPC_ENC_MSG_IN_38_MSG_IN_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_38_MSG_IN_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_38_MSG_IN_BIT_OFFSET = 0;
  localparam int LDPC_ENC_MSG_IN_39_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_MSG_IN_39_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_MSG_IN_39_BYTE_OFFSET = 13'h009c;
  localparam int LDPC_ENC_MSG_IN_39_MSG_IN_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_MSG_IN_39_MSG_IN_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_MSG_IN_39_MSG_IN_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_0_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_0_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_0_BYTE_OFFSET = 13'h00a0;
  localparam int LDPC_ENC_CODEWRD_OUT_0_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_0_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_0_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_1_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_1_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_1_BYTE_OFFSET = 13'h00a4;
  localparam int LDPC_ENC_CODEWRD_OUT_1_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_1_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_1_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_2_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_2_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_2_BYTE_OFFSET = 13'h00a8;
  localparam int LDPC_ENC_CODEWRD_OUT_2_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_2_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_2_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_3_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_3_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_3_BYTE_OFFSET = 13'h00ac;
  localparam int LDPC_ENC_CODEWRD_OUT_3_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_3_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_3_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_4_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_4_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_4_BYTE_OFFSET = 13'h00b0;
  localparam int LDPC_ENC_CODEWRD_OUT_4_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_4_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_4_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_5_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_5_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_5_BYTE_OFFSET = 13'h00b4;
  localparam int LDPC_ENC_CODEWRD_OUT_5_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_5_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_5_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_6_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_6_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_6_BYTE_OFFSET = 13'h00b8;
  localparam int LDPC_ENC_CODEWRD_OUT_6_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_6_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_6_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_7_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_7_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_7_BYTE_OFFSET = 13'h00bc;
  localparam int LDPC_ENC_CODEWRD_OUT_7_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_7_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_7_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_8_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_8_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_8_BYTE_OFFSET = 13'h00c0;
  localparam int LDPC_ENC_CODEWRD_OUT_8_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_8_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_8_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_9_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_9_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_9_BYTE_OFFSET = 13'h00c4;
  localparam int LDPC_ENC_CODEWRD_OUT_9_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_9_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_9_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_10_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_10_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_10_BYTE_OFFSET = 13'h00c8;
  localparam int LDPC_ENC_CODEWRD_OUT_10_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_10_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_10_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_11_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_11_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_11_BYTE_OFFSET = 13'h00cc;
  localparam int LDPC_ENC_CODEWRD_OUT_11_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_11_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_11_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_12_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_12_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_12_BYTE_OFFSET = 13'h00d0;
  localparam int LDPC_ENC_CODEWRD_OUT_12_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_12_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_12_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_13_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_13_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_13_BYTE_OFFSET = 13'h00d4;
  localparam int LDPC_ENC_CODEWRD_OUT_13_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_13_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_13_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_14_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_14_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_14_BYTE_OFFSET = 13'h00d8;
  localparam int LDPC_ENC_CODEWRD_OUT_14_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_14_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_14_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_15_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_15_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_15_BYTE_OFFSET = 13'h00dc;
  localparam int LDPC_ENC_CODEWRD_OUT_15_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_15_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_15_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_16_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_16_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_16_BYTE_OFFSET = 13'h00e0;
  localparam int LDPC_ENC_CODEWRD_OUT_16_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_16_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_16_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_17_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_17_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_17_BYTE_OFFSET = 13'h00e4;
  localparam int LDPC_ENC_CODEWRD_OUT_17_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_17_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_17_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_18_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_18_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_18_BYTE_OFFSET = 13'h00e8;
  localparam int LDPC_ENC_CODEWRD_OUT_18_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_18_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_18_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_19_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_19_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_19_BYTE_OFFSET = 13'h00ec;
  localparam int LDPC_ENC_CODEWRD_OUT_19_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_19_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_19_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_20_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_20_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_20_BYTE_OFFSET = 13'h00f0;
  localparam int LDPC_ENC_CODEWRD_OUT_20_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_20_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_20_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_21_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_21_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_21_BYTE_OFFSET = 13'h00f4;
  localparam int LDPC_ENC_CODEWRD_OUT_21_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_21_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_21_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_22_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_22_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_22_BYTE_OFFSET = 13'h00f8;
  localparam int LDPC_ENC_CODEWRD_OUT_22_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_22_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_22_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_23_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_23_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_23_BYTE_OFFSET = 13'h00fc;
  localparam int LDPC_ENC_CODEWRD_OUT_23_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_23_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_23_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_24_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_24_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_24_BYTE_OFFSET = 13'h0100;
  localparam int LDPC_ENC_CODEWRD_OUT_24_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_24_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_24_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_25_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_25_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_25_BYTE_OFFSET = 13'h0104;
  localparam int LDPC_ENC_CODEWRD_OUT_25_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_25_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_25_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_26_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_26_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_26_BYTE_OFFSET = 13'h0108;
  localparam int LDPC_ENC_CODEWRD_OUT_26_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_26_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_26_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_27_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_27_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_27_BYTE_OFFSET = 13'h010c;
  localparam int LDPC_ENC_CODEWRD_OUT_27_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_27_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_27_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_28_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_28_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_28_BYTE_OFFSET = 13'h0110;
  localparam int LDPC_ENC_CODEWRD_OUT_28_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_28_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_28_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_29_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_29_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_29_BYTE_OFFSET = 13'h0114;
  localparam int LDPC_ENC_CODEWRD_OUT_29_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_29_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_29_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_30_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_30_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_30_BYTE_OFFSET = 13'h0118;
  localparam int LDPC_ENC_CODEWRD_OUT_30_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_30_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_30_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_31_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_31_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_31_BYTE_OFFSET = 13'h011c;
  localparam int LDPC_ENC_CODEWRD_OUT_31_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_31_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_31_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_32_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_32_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_32_BYTE_OFFSET = 13'h0120;
  localparam int LDPC_ENC_CODEWRD_OUT_32_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_32_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_32_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_33_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_33_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_33_BYTE_OFFSET = 13'h0124;
  localparam int LDPC_ENC_CODEWRD_OUT_33_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_33_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_33_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_34_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_34_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_34_BYTE_OFFSET = 13'h0128;
  localparam int LDPC_ENC_CODEWRD_OUT_34_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_34_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_34_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_35_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_35_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_35_BYTE_OFFSET = 13'h012c;
  localparam int LDPC_ENC_CODEWRD_OUT_35_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_35_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_35_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_36_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_36_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_36_BYTE_OFFSET = 13'h0130;
  localparam int LDPC_ENC_CODEWRD_OUT_36_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_36_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_36_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_37_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_37_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_37_BYTE_OFFSET = 13'h0134;
  localparam int LDPC_ENC_CODEWRD_OUT_37_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_37_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_37_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_38_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_38_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_38_BYTE_OFFSET = 13'h0138;
  localparam int LDPC_ENC_CODEWRD_OUT_38_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_38_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_38_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_39_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_39_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_39_BYTE_OFFSET = 13'h013c;
  localparam int LDPC_ENC_CODEWRD_OUT_39_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_39_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_39_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_40_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_40_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_40_BYTE_OFFSET = 13'h0140;
  localparam int LDPC_ENC_CODEWRD_OUT_40_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_40_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_40_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_41_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_41_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_41_BYTE_OFFSET = 13'h0144;
  localparam int LDPC_ENC_CODEWRD_OUT_41_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_41_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_41_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_42_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_42_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_42_BYTE_OFFSET = 13'h0148;
  localparam int LDPC_ENC_CODEWRD_OUT_42_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_42_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_42_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_43_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_43_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_43_BYTE_OFFSET = 13'h014c;
  localparam int LDPC_ENC_CODEWRD_OUT_43_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_43_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_43_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_44_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_44_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_44_BYTE_OFFSET = 13'h0150;
  localparam int LDPC_ENC_CODEWRD_OUT_44_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_44_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_44_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_45_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_45_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_45_BYTE_OFFSET = 13'h0154;
  localparam int LDPC_ENC_CODEWRD_OUT_45_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_45_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_45_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_46_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_46_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_46_BYTE_OFFSET = 13'h0158;
  localparam int LDPC_ENC_CODEWRD_OUT_46_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_46_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_46_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_47_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_47_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_47_BYTE_OFFSET = 13'h015c;
  localparam int LDPC_ENC_CODEWRD_OUT_47_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_47_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_47_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_48_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_48_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_48_BYTE_OFFSET = 13'h0160;
  localparam int LDPC_ENC_CODEWRD_OUT_48_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_48_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_48_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_49_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_49_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_49_BYTE_OFFSET = 13'h0164;
  localparam int LDPC_ENC_CODEWRD_OUT_49_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_49_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_49_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_50_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_50_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_50_BYTE_OFFSET = 13'h0168;
  localparam int LDPC_ENC_CODEWRD_OUT_50_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_50_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_50_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_51_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_51_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_51_BYTE_OFFSET = 13'h016c;
  localparam int LDPC_ENC_CODEWRD_OUT_51_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_51_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_51_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_52_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_52_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_52_BYTE_OFFSET = 13'h0170;
  localparam int LDPC_ENC_CODEWRD_OUT_52_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_52_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_52_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_53_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_53_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_53_BYTE_OFFSET = 13'h0174;
  localparam int LDPC_ENC_CODEWRD_OUT_53_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_53_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_53_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_54_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_54_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_54_BYTE_OFFSET = 13'h0178;
  localparam int LDPC_ENC_CODEWRD_OUT_54_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_54_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_54_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_55_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_55_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_55_BYTE_OFFSET = 13'h017c;
  localparam int LDPC_ENC_CODEWRD_OUT_55_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_55_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_55_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_56_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_56_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_56_BYTE_OFFSET = 13'h0180;
  localparam int LDPC_ENC_CODEWRD_OUT_56_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_56_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_56_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_57_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_57_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_57_BYTE_OFFSET = 13'h0184;
  localparam int LDPC_ENC_CODEWRD_OUT_57_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_57_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_57_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_58_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_58_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_58_BYTE_OFFSET = 13'h0188;
  localparam int LDPC_ENC_CODEWRD_OUT_58_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_58_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_58_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_59_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_59_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_59_BYTE_OFFSET = 13'h018c;
  localparam int LDPC_ENC_CODEWRD_OUT_59_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_59_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_59_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_60_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_60_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_60_BYTE_OFFSET = 13'h0190;
  localparam int LDPC_ENC_CODEWRD_OUT_60_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_60_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_60_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_61_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_61_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_61_BYTE_OFFSET = 13'h0194;
  localparam int LDPC_ENC_CODEWRD_OUT_61_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_61_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_61_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_62_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_62_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_62_BYTE_OFFSET = 13'h0198;
  localparam int LDPC_ENC_CODEWRD_OUT_62_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_62_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_62_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_63_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_63_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_63_BYTE_OFFSET = 13'h019c;
  localparam int LDPC_ENC_CODEWRD_OUT_63_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_63_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_63_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_64_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_64_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_64_BYTE_OFFSET = 13'h01a0;
  localparam int LDPC_ENC_CODEWRD_OUT_64_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_64_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_64_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_65_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_65_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_65_BYTE_OFFSET = 13'h01a4;
  localparam int LDPC_ENC_CODEWRD_OUT_65_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_65_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_65_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_66_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_66_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_66_BYTE_OFFSET = 13'h01a8;
  localparam int LDPC_ENC_CODEWRD_OUT_66_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_66_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_66_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_67_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_67_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_67_BYTE_OFFSET = 13'h01ac;
  localparam int LDPC_ENC_CODEWRD_OUT_67_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_67_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_67_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_68_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_68_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_68_BYTE_OFFSET = 13'h01b0;
  localparam int LDPC_ENC_CODEWRD_OUT_68_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_68_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_68_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_69_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_69_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_69_BYTE_OFFSET = 13'h01b4;
  localparam int LDPC_ENC_CODEWRD_OUT_69_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_69_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_69_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_70_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_70_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_70_BYTE_OFFSET = 13'h01b8;
  localparam int LDPC_ENC_CODEWRD_OUT_70_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_70_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_70_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_71_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_71_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_71_BYTE_OFFSET = 13'h01bc;
  localparam int LDPC_ENC_CODEWRD_OUT_71_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_71_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_71_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_72_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_72_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_72_BYTE_OFFSET = 13'h01c0;
  localparam int LDPC_ENC_CODEWRD_OUT_72_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_72_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_72_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_73_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_73_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_73_BYTE_OFFSET = 13'h01c4;
  localparam int LDPC_ENC_CODEWRD_OUT_73_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_73_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_73_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_74_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_74_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_74_BYTE_OFFSET = 13'h01c8;
  localparam int LDPC_ENC_CODEWRD_OUT_74_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_74_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_74_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_75_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_75_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_75_BYTE_OFFSET = 13'h01cc;
  localparam int LDPC_ENC_CODEWRD_OUT_75_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_75_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_75_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_76_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_76_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_76_BYTE_OFFSET = 13'h01d0;
  localparam int LDPC_ENC_CODEWRD_OUT_76_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_76_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_76_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_77_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_77_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_77_BYTE_OFFSET = 13'h01d4;
  localparam int LDPC_ENC_CODEWRD_OUT_77_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_77_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_77_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_78_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_78_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_78_BYTE_OFFSET = 13'h01d8;
  localparam int LDPC_ENC_CODEWRD_OUT_78_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_78_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_78_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_79_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_79_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_79_BYTE_OFFSET = 13'h01dc;
  localparam int LDPC_ENC_CODEWRD_OUT_79_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_79_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_79_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_80_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_80_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_80_BYTE_OFFSET = 13'h01e0;
  localparam int LDPC_ENC_CODEWRD_OUT_80_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_80_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_80_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_81_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_81_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_81_BYTE_OFFSET = 13'h01e4;
  localparam int LDPC_ENC_CODEWRD_OUT_81_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_81_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_81_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_82_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_82_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_82_BYTE_OFFSET = 13'h01e8;
  localparam int LDPC_ENC_CODEWRD_OUT_82_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_82_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_82_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_83_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_83_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_83_BYTE_OFFSET = 13'h01ec;
  localparam int LDPC_ENC_CODEWRD_OUT_83_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_83_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_83_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_84_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_84_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_84_BYTE_OFFSET = 13'h01f0;
  localparam int LDPC_ENC_CODEWRD_OUT_84_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_84_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_84_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_85_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_85_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_85_BYTE_OFFSET = 13'h01f4;
  localparam int LDPC_ENC_CODEWRD_OUT_85_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_85_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_85_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_86_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_86_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_86_BYTE_OFFSET = 13'h01f8;
  localparam int LDPC_ENC_CODEWRD_OUT_86_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_86_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_86_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_87_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_87_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_87_BYTE_OFFSET = 13'h01fc;
  localparam int LDPC_ENC_CODEWRD_OUT_87_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_87_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_87_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_88_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_88_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_88_BYTE_OFFSET = 13'h0200;
  localparam int LDPC_ENC_CODEWRD_OUT_88_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_88_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_88_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_89_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_89_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_89_BYTE_OFFSET = 13'h0204;
  localparam int LDPC_ENC_CODEWRD_OUT_89_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_89_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_89_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_90_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_90_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_90_BYTE_OFFSET = 13'h0208;
  localparam int LDPC_ENC_CODEWRD_OUT_90_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_90_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_90_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_91_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_91_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_91_BYTE_OFFSET = 13'h020c;
  localparam int LDPC_ENC_CODEWRD_OUT_91_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_91_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_91_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_92_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_92_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_92_BYTE_OFFSET = 13'h0210;
  localparam int LDPC_ENC_CODEWRD_OUT_92_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_92_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_92_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_93_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_93_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_93_BYTE_OFFSET = 13'h0214;
  localparam int LDPC_ENC_CODEWRD_OUT_93_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_93_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_93_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_94_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_94_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_94_BYTE_OFFSET = 13'h0218;
  localparam int LDPC_ENC_CODEWRD_OUT_94_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_94_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_94_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_95_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_95_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_95_BYTE_OFFSET = 13'h021c;
  localparam int LDPC_ENC_CODEWRD_OUT_95_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_95_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_95_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_96_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_96_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_96_BYTE_OFFSET = 13'h0220;
  localparam int LDPC_ENC_CODEWRD_OUT_96_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_96_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_96_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_97_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_97_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_97_BYTE_OFFSET = 13'h0224;
  localparam int LDPC_ENC_CODEWRD_OUT_97_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_97_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_97_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_98_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_98_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_98_BYTE_OFFSET = 13'h0228;
  localparam int LDPC_ENC_CODEWRD_OUT_98_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_98_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_98_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_99_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_99_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_99_BYTE_OFFSET = 13'h022c;
  localparam int LDPC_ENC_CODEWRD_OUT_99_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_99_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_99_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_100_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_100_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_100_BYTE_OFFSET = 13'h0230;
  localparam int LDPC_ENC_CODEWRD_OUT_100_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_100_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_100_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_101_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_101_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_101_BYTE_OFFSET = 13'h0234;
  localparam int LDPC_ENC_CODEWRD_OUT_101_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_101_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_101_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_102_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_102_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_102_BYTE_OFFSET = 13'h0238;
  localparam int LDPC_ENC_CODEWRD_OUT_102_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_102_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_102_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_103_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_103_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_103_BYTE_OFFSET = 13'h023c;
  localparam int LDPC_ENC_CODEWRD_OUT_103_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_103_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_103_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_104_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_104_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_104_BYTE_OFFSET = 13'h0240;
  localparam int LDPC_ENC_CODEWRD_OUT_104_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_104_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_104_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_105_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_105_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_105_BYTE_OFFSET = 13'h0244;
  localparam int LDPC_ENC_CODEWRD_OUT_105_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_105_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_105_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_106_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_106_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_106_BYTE_OFFSET = 13'h0248;
  localparam int LDPC_ENC_CODEWRD_OUT_106_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_106_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_106_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_107_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_107_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_107_BYTE_OFFSET = 13'h024c;
  localparam int LDPC_ENC_CODEWRD_OUT_107_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_107_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_107_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_108_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_108_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_108_BYTE_OFFSET = 13'h0250;
  localparam int LDPC_ENC_CODEWRD_OUT_108_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_108_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_108_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_109_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_109_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_109_BYTE_OFFSET = 13'h0254;
  localparam int LDPC_ENC_CODEWRD_OUT_109_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_109_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_109_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_110_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_110_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_110_BYTE_OFFSET = 13'h0258;
  localparam int LDPC_ENC_CODEWRD_OUT_110_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_110_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_110_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_111_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_111_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_111_BYTE_OFFSET = 13'h025c;
  localparam int LDPC_ENC_CODEWRD_OUT_111_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_111_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_111_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_112_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_112_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_112_BYTE_OFFSET = 13'h0260;
  localparam int LDPC_ENC_CODEWRD_OUT_112_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_112_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_112_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_113_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_113_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_113_BYTE_OFFSET = 13'h0264;
  localparam int LDPC_ENC_CODEWRD_OUT_113_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_113_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_113_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_114_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_114_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_114_BYTE_OFFSET = 13'h0268;
  localparam int LDPC_ENC_CODEWRD_OUT_114_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_114_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_114_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_115_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_115_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_115_BYTE_OFFSET = 13'h026c;
  localparam int LDPC_ENC_CODEWRD_OUT_115_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_115_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_115_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_116_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_116_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_116_BYTE_OFFSET = 13'h0270;
  localparam int LDPC_ENC_CODEWRD_OUT_116_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_116_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_116_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_117_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_117_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_117_BYTE_OFFSET = 13'h0274;
  localparam int LDPC_ENC_CODEWRD_OUT_117_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_117_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_117_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_118_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_118_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_118_BYTE_OFFSET = 13'h0278;
  localparam int LDPC_ENC_CODEWRD_OUT_118_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_118_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_118_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_119_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_119_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_119_BYTE_OFFSET = 13'h027c;
  localparam int LDPC_ENC_CODEWRD_OUT_119_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_119_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_119_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_120_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_120_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_120_BYTE_OFFSET = 13'h0280;
  localparam int LDPC_ENC_CODEWRD_OUT_120_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_120_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_120_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_121_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_121_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_121_BYTE_OFFSET = 13'h0284;
  localparam int LDPC_ENC_CODEWRD_OUT_121_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_121_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_121_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_122_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_122_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_122_BYTE_OFFSET = 13'h0288;
  localparam int LDPC_ENC_CODEWRD_OUT_122_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_122_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_122_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_123_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_123_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_123_BYTE_OFFSET = 13'h028c;
  localparam int LDPC_ENC_CODEWRD_OUT_123_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_123_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_123_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_124_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_124_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_124_BYTE_OFFSET = 13'h0290;
  localparam int LDPC_ENC_CODEWRD_OUT_124_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_124_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_124_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_125_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_125_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_125_BYTE_OFFSET = 13'h0294;
  localparam int LDPC_ENC_CODEWRD_OUT_125_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_125_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_125_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_126_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_126_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_126_BYTE_OFFSET = 13'h0298;
  localparam int LDPC_ENC_CODEWRD_OUT_126_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_126_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_126_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_127_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_127_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_127_BYTE_OFFSET = 13'h029c;
  localparam int LDPC_ENC_CODEWRD_OUT_127_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_127_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_127_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_128_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_128_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_128_BYTE_OFFSET = 13'h02a0;
  localparam int LDPC_ENC_CODEWRD_OUT_128_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_128_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_128_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_129_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_129_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_129_BYTE_OFFSET = 13'h02a4;
  localparam int LDPC_ENC_CODEWRD_OUT_129_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_129_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_129_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_130_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_130_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_130_BYTE_OFFSET = 13'h02a8;
  localparam int LDPC_ENC_CODEWRD_OUT_130_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_130_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_130_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_131_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_131_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_131_BYTE_OFFSET = 13'h02ac;
  localparam int LDPC_ENC_CODEWRD_OUT_131_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_131_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_131_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_132_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_132_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_132_BYTE_OFFSET = 13'h02b0;
  localparam int LDPC_ENC_CODEWRD_OUT_132_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_132_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_132_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_133_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_133_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_133_BYTE_OFFSET = 13'h02b4;
  localparam int LDPC_ENC_CODEWRD_OUT_133_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_133_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_133_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_134_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_134_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_134_BYTE_OFFSET = 13'h02b8;
  localparam int LDPC_ENC_CODEWRD_OUT_134_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_134_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_134_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_135_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_135_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_135_BYTE_OFFSET = 13'h02bc;
  localparam int LDPC_ENC_CODEWRD_OUT_135_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_135_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_135_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_136_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_136_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_136_BYTE_OFFSET = 13'h02c0;
  localparam int LDPC_ENC_CODEWRD_OUT_136_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_136_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_136_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_137_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_137_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_137_BYTE_OFFSET = 13'h02c4;
  localparam int LDPC_ENC_CODEWRD_OUT_137_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_137_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_137_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_138_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_138_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_138_BYTE_OFFSET = 13'h02c8;
  localparam int LDPC_ENC_CODEWRD_OUT_138_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_138_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_138_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_139_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_139_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_139_BYTE_OFFSET = 13'h02cc;
  localparam int LDPC_ENC_CODEWRD_OUT_139_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_139_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_139_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_140_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_140_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_140_BYTE_OFFSET = 13'h02d0;
  localparam int LDPC_ENC_CODEWRD_OUT_140_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_140_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_140_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_141_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_141_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_141_BYTE_OFFSET = 13'h02d4;
  localparam int LDPC_ENC_CODEWRD_OUT_141_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_141_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_141_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_142_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_142_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_142_BYTE_OFFSET = 13'h02d8;
  localparam int LDPC_ENC_CODEWRD_OUT_142_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_142_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_142_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_143_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_143_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_143_BYTE_OFFSET = 13'h02dc;
  localparam int LDPC_ENC_CODEWRD_OUT_143_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_143_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_143_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_144_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_144_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_144_BYTE_OFFSET = 13'h02e0;
  localparam int LDPC_ENC_CODEWRD_OUT_144_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_144_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_144_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_145_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_145_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_145_BYTE_OFFSET = 13'h02e4;
  localparam int LDPC_ENC_CODEWRD_OUT_145_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_145_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_145_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_146_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_146_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_146_BYTE_OFFSET = 13'h02e8;
  localparam int LDPC_ENC_CODEWRD_OUT_146_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_146_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_146_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_147_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_147_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_147_BYTE_OFFSET = 13'h02ec;
  localparam int LDPC_ENC_CODEWRD_OUT_147_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_147_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_147_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_148_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_148_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_148_BYTE_OFFSET = 13'h02f0;
  localparam int LDPC_ENC_CODEWRD_OUT_148_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_148_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_148_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_149_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_149_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_149_BYTE_OFFSET = 13'h02f4;
  localparam int LDPC_ENC_CODEWRD_OUT_149_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_149_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_149_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_150_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_150_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_150_BYTE_OFFSET = 13'h02f8;
  localparam int LDPC_ENC_CODEWRD_OUT_150_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_150_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_150_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_151_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_151_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_151_BYTE_OFFSET = 13'h02fc;
  localparam int LDPC_ENC_CODEWRD_OUT_151_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_151_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_151_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_152_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_152_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_152_BYTE_OFFSET = 13'h0300;
  localparam int LDPC_ENC_CODEWRD_OUT_152_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_152_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_152_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_153_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_153_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_153_BYTE_OFFSET = 13'h0304;
  localparam int LDPC_ENC_CODEWRD_OUT_153_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_153_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_153_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_154_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_154_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_154_BYTE_OFFSET = 13'h0308;
  localparam int LDPC_ENC_CODEWRD_OUT_154_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_154_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_154_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_155_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_155_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_155_BYTE_OFFSET = 13'h030c;
  localparam int LDPC_ENC_CODEWRD_OUT_155_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_155_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_155_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_156_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_156_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_156_BYTE_OFFSET = 13'h0310;
  localparam int LDPC_ENC_CODEWRD_OUT_156_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_156_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_156_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_157_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_157_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_157_BYTE_OFFSET = 13'h0314;
  localparam int LDPC_ENC_CODEWRD_OUT_157_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_157_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_157_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_158_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_158_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_158_BYTE_OFFSET = 13'h0318;
  localparam int LDPC_ENC_CODEWRD_OUT_158_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_158_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_158_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_159_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_159_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_159_BYTE_OFFSET = 13'h031c;
  localparam int LDPC_ENC_CODEWRD_OUT_159_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_159_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_159_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_160_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_160_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_160_BYTE_OFFSET = 13'h0320;
  localparam int LDPC_ENC_CODEWRD_OUT_160_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_160_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_160_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_161_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_161_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_161_BYTE_OFFSET = 13'h0324;
  localparam int LDPC_ENC_CODEWRD_OUT_161_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_161_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_161_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_162_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_162_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_162_BYTE_OFFSET = 13'h0328;
  localparam int LDPC_ENC_CODEWRD_OUT_162_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_162_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_162_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_163_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_163_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_163_BYTE_OFFSET = 13'h032c;
  localparam int LDPC_ENC_CODEWRD_OUT_163_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_163_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_163_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_164_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_164_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_164_BYTE_OFFSET = 13'h0330;
  localparam int LDPC_ENC_CODEWRD_OUT_164_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_164_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_164_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_165_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_165_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_165_BYTE_OFFSET = 13'h0334;
  localparam int LDPC_ENC_CODEWRD_OUT_165_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_165_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_165_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_166_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_166_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_166_BYTE_OFFSET = 13'h0338;
  localparam int LDPC_ENC_CODEWRD_OUT_166_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_166_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_166_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_167_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_167_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_167_BYTE_OFFSET = 13'h033c;
  localparam int LDPC_ENC_CODEWRD_OUT_167_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_167_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_167_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_168_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_168_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_168_BYTE_OFFSET = 13'h0340;
  localparam int LDPC_ENC_CODEWRD_OUT_168_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_168_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_168_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_169_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_169_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_169_BYTE_OFFSET = 13'h0344;
  localparam int LDPC_ENC_CODEWRD_OUT_169_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_169_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_169_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_170_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_170_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_170_BYTE_OFFSET = 13'h0348;
  localparam int LDPC_ENC_CODEWRD_OUT_170_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_170_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_170_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_171_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_171_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_171_BYTE_OFFSET = 13'h034c;
  localparam int LDPC_ENC_CODEWRD_OUT_171_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_171_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_171_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_172_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_172_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_172_BYTE_OFFSET = 13'h0350;
  localparam int LDPC_ENC_CODEWRD_OUT_172_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_172_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_172_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_173_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_173_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_173_BYTE_OFFSET = 13'h0354;
  localparam int LDPC_ENC_CODEWRD_OUT_173_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_173_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_173_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_174_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_174_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_174_BYTE_OFFSET = 13'h0358;
  localparam int LDPC_ENC_CODEWRD_OUT_174_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_174_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_174_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_175_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_175_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_175_BYTE_OFFSET = 13'h035c;
  localparam int LDPC_ENC_CODEWRD_OUT_175_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_175_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_175_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_176_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_176_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_176_BYTE_OFFSET = 13'h0360;
  localparam int LDPC_ENC_CODEWRD_OUT_176_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_176_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_176_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_177_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_177_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_177_BYTE_OFFSET = 13'h0364;
  localparam int LDPC_ENC_CODEWRD_OUT_177_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_177_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_177_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_178_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_178_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_178_BYTE_OFFSET = 13'h0368;
  localparam int LDPC_ENC_CODEWRD_OUT_178_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_178_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_178_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_179_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_179_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_179_BYTE_OFFSET = 13'h036c;
  localparam int LDPC_ENC_CODEWRD_OUT_179_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_179_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_179_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_180_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_180_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_180_BYTE_OFFSET = 13'h0370;
  localparam int LDPC_ENC_CODEWRD_OUT_180_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_180_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_180_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_181_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_181_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_181_BYTE_OFFSET = 13'h0374;
  localparam int LDPC_ENC_CODEWRD_OUT_181_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_181_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_181_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_182_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_182_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_182_BYTE_OFFSET = 13'h0378;
  localparam int LDPC_ENC_CODEWRD_OUT_182_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_182_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_182_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_183_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_183_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_183_BYTE_OFFSET = 13'h037c;
  localparam int LDPC_ENC_CODEWRD_OUT_183_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_183_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_183_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_184_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_184_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_184_BYTE_OFFSET = 13'h0380;
  localparam int LDPC_ENC_CODEWRD_OUT_184_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_184_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_184_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_185_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_185_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_185_BYTE_OFFSET = 13'h0384;
  localparam int LDPC_ENC_CODEWRD_OUT_185_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_185_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_185_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_186_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_186_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_186_BYTE_OFFSET = 13'h0388;
  localparam int LDPC_ENC_CODEWRD_OUT_186_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_186_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_186_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_187_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_187_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_187_BYTE_OFFSET = 13'h038c;
  localparam int LDPC_ENC_CODEWRD_OUT_187_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_187_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_187_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_188_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_188_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_188_BYTE_OFFSET = 13'h0390;
  localparam int LDPC_ENC_CODEWRD_OUT_188_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_188_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_188_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_189_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_189_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_189_BYTE_OFFSET = 13'h0394;
  localparam int LDPC_ENC_CODEWRD_OUT_189_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_189_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_189_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_190_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_190_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_190_BYTE_OFFSET = 13'h0398;
  localparam int LDPC_ENC_CODEWRD_OUT_190_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_190_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_190_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_191_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_191_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_191_BYTE_OFFSET = 13'h039c;
  localparam int LDPC_ENC_CODEWRD_OUT_191_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_191_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_191_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_192_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_192_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_192_BYTE_OFFSET = 13'h03a0;
  localparam int LDPC_ENC_CODEWRD_OUT_192_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_192_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_192_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_193_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_193_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_193_BYTE_OFFSET = 13'h03a4;
  localparam int LDPC_ENC_CODEWRD_OUT_193_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_193_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_193_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_194_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_194_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_194_BYTE_OFFSET = 13'h03a8;
  localparam int LDPC_ENC_CODEWRD_OUT_194_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_194_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_194_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_195_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_195_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_195_BYTE_OFFSET = 13'h03ac;
  localparam int LDPC_ENC_CODEWRD_OUT_195_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_195_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_195_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_196_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_196_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_196_BYTE_OFFSET = 13'h03b0;
  localparam int LDPC_ENC_CODEWRD_OUT_196_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_196_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_196_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_197_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_197_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_197_BYTE_OFFSET = 13'h03b4;
  localparam int LDPC_ENC_CODEWRD_OUT_197_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_197_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_197_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_198_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_198_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_198_BYTE_OFFSET = 13'h03b8;
  localparam int LDPC_ENC_CODEWRD_OUT_198_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_198_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_198_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_199_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_199_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_199_BYTE_OFFSET = 13'h03bc;
  localparam int LDPC_ENC_CODEWRD_OUT_199_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_199_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_199_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_200_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_200_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_200_BYTE_OFFSET = 13'h03c0;
  localparam int LDPC_ENC_CODEWRD_OUT_200_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_200_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_200_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_201_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_201_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_201_BYTE_OFFSET = 13'h03c4;
  localparam int LDPC_ENC_CODEWRD_OUT_201_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_201_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_201_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_202_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_202_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_202_BYTE_OFFSET = 13'h03c8;
  localparam int LDPC_ENC_CODEWRD_OUT_202_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_202_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_202_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_203_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_203_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_203_BYTE_OFFSET = 13'h03cc;
  localparam int LDPC_ENC_CODEWRD_OUT_203_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_203_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_203_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_204_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_204_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_204_BYTE_OFFSET = 13'h03d0;
  localparam int LDPC_ENC_CODEWRD_OUT_204_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_204_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_204_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_205_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_205_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_205_BYTE_OFFSET = 13'h03d4;
  localparam int LDPC_ENC_CODEWRD_OUT_205_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_205_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_205_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_206_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_206_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_206_BYTE_OFFSET = 13'h03d8;
  localparam int LDPC_ENC_CODEWRD_OUT_206_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_206_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_206_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_OUT_207_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_OUT_207_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_OUT_207_BYTE_OFFSET = 13'h03dc;
  localparam int LDPC_ENC_CODEWRD_OUT_207_ENC_CODEWORD_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_OUT_207_ENC_CODEWORD_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_OUT_207_ENC_CODEWORD_BIT_OFFSET = 0;
  localparam int LDPC_ENC_CODEWRD_VLD_BYTE_WIDTH = 4;
  localparam int LDPC_ENC_CODEWRD_VLD_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_ENC_CODEWRD_VLD_BYTE_OFFSET = 13'h03e0;
  localparam int LDPC_ENC_CODEWRD_VLD_ENC_CODEWORD_VALID_BIT_WIDTH = 1;
  localparam bit LDPC_ENC_CODEWRD_VLD_ENC_CODEWORD_VALID_BIT_MASK = 1'h1;
  localparam int LDPC_ENC_CODEWRD_VLD_ENC_CODEWORD_VALID_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_INTRODUCED_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_INTRODUCED_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_INTRODUCED_BYTE_OFFSET = 13'h03e4;
  localparam int LDPC_DEC_ERR_INTRODUCED_ERR_INTRO_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_INTRODUCED_ERR_INTRO_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_INTRODUCED_ERR_INTRO_BIT_OFFSET = 0;
  localparam int LDPC_DEC_SEL_FRMC_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_SEL_FRMC_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_SEL_FRMC_BYTE_OFFSET = 13'h03e8;
  localparam int LDPC_DEC_SEL_FRMC_SEL_Q0_FRMC_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_SEL_FRMC_SEL_Q0_FRMC_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_SEL_FRMC_SEL_Q0_FRMC_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_0_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_0_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_0_BYTE_OFFSET = 13'h03ec;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_0_ERR_INTRO_Q0_0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_0_ERR_INTRO_Q0_0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_0_ERR_INTRO_Q0_0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_1_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_1_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_1_BYTE_OFFSET = 13'h03f0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_1_ERR_INTRO_Q0_0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_1_ERR_INTRO_Q0_0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_1_ERR_INTRO_Q0_0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_2_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_2_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_2_BYTE_OFFSET = 13'h03f4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_2_ERR_INTRO_Q0_0_2_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_2_ERR_INTRO_Q0_0_2_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_2_ERR_INTRO_Q0_0_2_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_3_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_3_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_3_BYTE_OFFSET = 13'h03f8;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_3_ERR_INTRO_Q0_0_3_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_3_ERR_INTRO_Q0_0_3_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_3_ERR_INTRO_Q0_0_3_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_4_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_4_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_4_BYTE_OFFSET = 13'h03fc;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_4_ERR_INTRO_Q0_0_4_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_4_ERR_INTRO_Q0_0_4_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_4_ERR_INTRO_Q0_0_4_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_5_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_5_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_5_BYTE_OFFSET = 13'h0400;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_5_ERR_INTRO_Q0_0_5_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_5_ERR_INTRO_Q0_0_5_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_5_ERR_INTRO_Q0_0_5_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_6_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_6_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_6_BYTE_OFFSET = 13'h0404;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_6_ERR_INTRO_Q0_0_6_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_6_ERR_INTRO_Q0_0_6_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_6_ERR_INTRO_Q0_0_6_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_7_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_7_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_7_BYTE_OFFSET = 13'h0408;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_7_ERR_INTRO_Q0_0_7_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_7_ERR_INTRO_Q0_0_7_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_7_ERR_INTRO_Q0_0_7_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_8_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_8_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_8_BYTE_OFFSET = 13'h040c;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_8_ERR_INTRO_Q0_0_8_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_8_ERR_INTRO_Q0_0_8_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_8_ERR_INTRO_Q0_0_8_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_9_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_9_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_9_BYTE_OFFSET = 13'h0410;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_9_ERR_INTRO_Q0_0_9_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_9_ERR_INTRO_Q0_0_9_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_9_ERR_INTRO_Q0_0_9_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_10_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_10_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_10_BYTE_OFFSET = 13'h0414;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_10_ERR_INTRO_Q0_0_10_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_10_ERR_INTRO_Q0_0_10_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_10_ERR_INTRO_Q0_0_10_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_11_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_11_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_11_BYTE_OFFSET = 13'h0418;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_11_ERR_INTRO_Q0_0_11_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_11_ERR_INTRO_Q0_0_11_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_11_ERR_INTRO_Q0_0_11_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_12_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_12_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_12_BYTE_OFFSET = 13'h041c;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_12_ERR_INTRO_Q0_0_12_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_12_ERR_INTRO_Q0_0_12_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_12_ERR_INTRO_Q0_0_12_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_13_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_13_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_13_BYTE_OFFSET = 13'h0420;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_13_ERR_INTRO_Q0_0_13_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_13_ERR_INTRO_Q0_0_13_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_13_ERR_INTRO_Q0_0_13_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_14_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_14_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_14_BYTE_OFFSET = 13'h0424;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_14_ERR_INTRO_Q0_0_14_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_14_ERR_INTRO_Q0_0_14_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_14_ERR_INTRO_Q0_0_14_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_15_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_15_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_15_BYTE_OFFSET = 13'h0428;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_15_ERR_INTRO_Q0_0_15_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_15_ERR_INTRO_Q0_0_15_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_15_ERR_INTRO_Q0_0_15_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_16_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_16_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_16_BYTE_OFFSET = 13'h042c;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_16_ERR_INTRO_Q0_0_16_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_16_ERR_INTRO_Q0_0_16_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_16_ERR_INTRO_Q0_0_16_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_17_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_17_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_17_BYTE_OFFSET = 13'h0430;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_17_ERR_INTRO_Q0_0_17_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_17_ERR_INTRO_Q0_0_17_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_17_ERR_INTRO_Q0_0_17_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_18_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_18_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_18_BYTE_OFFSET = 13'h0434;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_18_ERR_INTRO_Q0_0_18_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_18_ERR_INTRO_Q0_0_18_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_18_ERR_INTRO_Q0_0_18_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_19_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_19_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_19_BYTE_OFFSET = 13'h0438;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_19_ERR_INTRO_Q0_0_19_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_19_ERR_INTRO_Q0_0_19_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_19_ERR_INTRO_Q0_0_19_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_20_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_20_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_20_BYTE_OFFSET = 13'h043c;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_20_ERR_INTRO_Q0_0_20_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_20_ERR_INTRO_Q0_0_20_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_20_ERR_INTRO_Q0_0_20_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_21_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_21_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_21_BYTE_OFFSET = 13'h0440;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_21_ERR_INTRO_Q0_0_21_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_21_ERR_INTRO_Q0_0_21_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_21_ERR_INTRO_Q0_0_21_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_22_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_22_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_22_BYTE_OFFSET = 13'h0444;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_22_ERR_INTRO_Q0_0_22_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_22_ERR_INTRO_Q0_0_22_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_22_ERR_INTRO_Q0_0_22_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_23_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_23_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_23_BYTE_OFFSET = 13'h0448;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_23_ERR_INTRO_Q0_0_23_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_23_ERR_INTRO_Q0_0_23_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_23_ERR_INTRO_Q0_0_23_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_24_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_24_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_24_BYTE_OFFSET = 13'h044c;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_24_ERR_INTRO_Q0_0_24_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_24_ERR_INTRO_Q0_0_24_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_24_ERR_INTRO_Q0_0_24_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_25_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_25_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_25_BYTE_OFFSET = 13'h0450;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_25_ERR_INTRO_Q0_0_25_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_25_ERR_INTRO_Q0_0_25_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_25_ERR_INTRO_Q0_0_25_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_26_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_26_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_26_BYTE_OFFSET = 13'h0454;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_26_ERR_INTRO_Q0_0_26_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_26_ERR_INTRO_Q0_0_26_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_26_ERR_INTRO_Q0_0_26_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_27_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_27_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_27_BYTE_OFFSET = 13'h0458;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_27_ERR_INTRO_Q0_0_27_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_27_ERR_INTRO_Q0_0_27_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_27_ERR_INTRO_Q0_0_27_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_28_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_28_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_28_BYTE_OFFSET = 13'h045c;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_28_ERR_INTRO_Q0_0_28_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_28_ERR_INTRO_Q0_0_28_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_28_ERR_INTRO_Q0_0_28_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_29_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_29_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_29_BYTE_OFFSET = 13'h0460;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_29_ERR_INTRO_Q0_0_29_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_29_ERR_INTRO_Q0_0_29_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_29_ERR_INTRO_Q0_0_29_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_30_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_30_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_30_BYTE_OFFSET = 13'h0464;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_30_ERR_INTRO_Q0_0_30_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_30_ERR_INTRO_Q0_0_30_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_30_ERR_INTRO_Q0_0_30_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_31_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_31_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_31_BYTE_OFFSET = 13'h0468;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_31_ERR_INTRO_Q0_0_31_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_31_ERR_INTRO_Q0_0_31_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_31_ERR_INTRO_Q0_0_31_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_32_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_32_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_32_BYTE_OFFSET = 13'h046c;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_32_ERR_INTRO_Q0_0_32_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_32_ERR_INTRO_Q0_0_32_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_32_ERR_INTRO_Q0_0_32_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_33_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_33_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_33_BYTE_OFFSET = 13'h0470;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_33_ERR_INTRO_Q0_0_33_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_33_ERR_INTRO_Q0_0_33_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_33_ERR_INTRO_Q0_0_33_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_34_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_34_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_34_BYTE_OFFSET = 13'h0474;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_34_ERR_INTRO_Q0_0_34_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_34_ERR_INTRO_Q0_0_34_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_34_ERR_INTRO_Q0_0_34_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_35_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_35_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_35_BYTE_OFFSET = 13'h0478;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_35_ERR_INTRO_Q0_0_35_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_35_ERR_INTRO_Q0_0_35_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_35_ERR_INTRO_Q0_0_35_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_36_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_36_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_36_BYTE_OFFSET = 13'h047c;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_36_ERR_INTRO_Q0_0_36_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_36_ERR_INTRO_Q0_0_36_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_36_ERR_INTRO_Q0_0_36_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_37_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_37_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_37_BYTE_OFFSET = 13'h0480;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_37_ERR_INTRO_Q0_0_37_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_37_ERR_INTRO_Q0_0_37_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_37_ERR_INTRO_Q0_0_37_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_38_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_38_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_38_BYTE_OFFSET = 13'h0484;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_38_ERR_INTRO_Q0_0_38_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_38_ERR_INTRO_Q0_0_38_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_38_ERR_INTRO_Q0_0_38_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_39_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_39_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_39_BYTE_OFFSET = 13'h0488;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_39_ERR_INTRO_Q0_0_39_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_39_ERR_INTRO_Q0_0_39_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_39_ERR_INTRO_Q0_0_39_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_40_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_40_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_40_BYTE_OFFSET = 13'h048c;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_40_ERR_INTRO_Q0_0_40_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_40_ERR_INTRO_Q0_0_40_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_40_ERR_INTRO_Q0_0_40_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_41_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_41_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_41_BYTE_OFFSET = 13'h0490;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_41_ERR_INTRO_Q0_0_41_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_41_ERR_INTRO_Q0_0_41_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_41_ERR_INTRO_Q0_0_41_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_42_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_42_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_42_BYTE_OFFSET = 13'h0494;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_42_ERR_INTRO_Q0_0_42_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_42_ERR_INTRO_Q0_0_42_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_42_ERR_INTRO_Q0_0_42_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_43_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_43_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_43_BYTE_OFFSET = 13'h0498;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_43_ERR_INTRO_Q0_0_43_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_43_ERR_INTRO_Q0_0_43_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_43_ERR_INTRO_Q0_0_43_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_44_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_44_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_44_BYTE_OFFSET = 13'h049c;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_44_ERR_INTRO_Q0_0_44_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_44_ERR_INTRO_Q0_0_44_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_44_ERR_INTRO_Q0_0_44_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_45_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_45_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_45_BYTE_OFFSET = 13'h04a0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_45_ERR_INTRO_Q0_0_45_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_45_ERR_INTRO_Q0_0_45_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_45_ERR_INTRO_Q0_0_45_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_46_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_46_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_46_BYTE_OFFSET = 13'h04a4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_46_ERR_INTRO_Q0_0_46_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_46_ERR_INTRO_Q0_0_46_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_46_ERR_INTRO_Q0_0_46_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_47_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_47_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_47_BYTE_OFFSET = 13'h04a8;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_47_ERR_INTRO_Q0_0_47_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_47_ERR_INTRO_Q0_0_47_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_47_ERR_INTRO_Q0_0_47_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_48_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_48_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_48_BYTE_OFFSET = 13'h04ac;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_48_ERR_INTRO_Q0_0_48_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_48_ERR_INTRO_Q0_0_48_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_48_ERR_INTRO_Q0_0_48_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_49_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_49_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_49_BYTE_OFFSET = 13'h04b0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_49_ERR_INTRO_Q0_0_49_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_49_ERR_INTRO_Q0_0_49_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_49_ERR_INTRO_Q0_0_49_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_50_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_50_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_50_BYTE_OFFSET = 13'h04b4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_50_ERR_INTRO_Q0_0_50_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_50_ERR_INTRO_Q0_0_50_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_50_ERR_INTRO_Q0_0_50_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_51_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_51_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_51_BYTE_OFFSET = 13'h04b8;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_51_ERR_INTRO_Q0_0_51_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_51_ERR_INTRO_Q0_0_51_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_51_ERR_INTRO_Q0_0_51_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_52_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_52_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_52_BYTE_OFFSET = 13'h04bc;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_52_ERR_INTRO_Q0_0_52_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_52_ERR_INTRO_Q0_0_52_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_52_ERR_INTRO_Q0_0_52_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_53_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_53_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_53_BYTE_OFFSET = 13'h04c0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_53_ERR_INTRO_Q0_0_53_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_53_ERR_INTRO_Q0_0_53_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_53_ERR_INTRO_Q0_0_53_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_54_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_54_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_54_BYTE_OFFSET = 13'h04c4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_54_ERR_INTRO_Q0_0_54_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_54_ERR_INTRO_Q0_0_54_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_54_ERR_INTRO_Q0_0_54_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_55_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_55_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_55_BYTE_OFFSET = 13'h04c8;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_55_ERR_INTRO_Q0_0_55_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_55_ERR_INTRO_Q0_0_55_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_55_ERR_INTRO_Q0_0_55_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_56_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_56_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_56_BYTE_OFFSET = 13'h04cc;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_56_ERR_INTRO_Q0_0_56_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_56_ERR_INTRO_Q0_0_56_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_56_ERR_INTRO_Q0_0_56_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_57_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_57_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_57_BYTE_OFFSET = 13'h04d0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_57_ERR_INTRO_Q0_0_57_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_57_ERR_INTRO_Q0_0_57_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_57_ERR_INTRO_Q0_0_57_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_58_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_58_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_58_BYTE_OFFSET = 13'h04d4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_58_ERR_INTRO_Q0_0_58_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_58_ERR_INTRO_Q0_0_58_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_58_ERR_INTRO_Q0_0_58_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_59_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_59_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_59_BYTE_OFFSET = 13'h04d8;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_59_ERR_INTRO_Q0_0_59_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_59_ERR_INTRO_Q0_0_59_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_59_ERR_INTRO_Q0_0_59_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_60_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_60_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_60_BYTE_OFFSET = 13'h04dc;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_60_ERR_INTRO_Q0_0_60_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_60_ERR_INTRO_Q0_0_60_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_60_ERR_INTRO_Q0_0_60_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_61_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_61_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_61_BYTE_OFFSET = 13'h04e0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_61_ERR_INTRO_Q0_0_61_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_61_ERR_INTRO_Q0_0_61_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_61_ERR_INTRO_Q0_0_61_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_62_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_62_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_62_BYTE_OFFSET = 13'h04e4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_62_ERR_INTRO_Q0_0_62_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_62_ERR_INTRO_Q0_0_62_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_62_ERR_INTRO_Q0_0_62_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_63_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_63_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_63_BYTE_OFFSET = 13'h04e8;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_63_ERR_INTRO_Q0_0_63_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_63_ERR_INTRO_Q0_0_63_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_63_ERR_INTRO_Q0_0_63_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_64_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_64_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_64_BYTE_OFFSET = 13'h04ec;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_64_ERR_INTRO_Q0_0_64_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_64_ERR_INTRO_Q0_0_64_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_64_ERR_INTRO_Q0_0_64_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_65_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_65_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_65_BYTE_OFFSET = 13'h04f0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_65_ERR_INTRO_Q0_0_65_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_65_ERR_INTRO_Q0_0_65_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_65_ERR_INTRO_Q0_0_65_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_66_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_66_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_66_BYTE_OFFSET = 13'h04f4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_66_ERR_INTRO_Q0_0_66_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_66_ERR_INTRO_Q0_0_66_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_66_ERR_INTRO_Q0_0_66_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_67_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_67_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_67_BYTE_OFFSET = 13'h04f8;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_67_ERR_INTRO_Q0_0_67_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_67_ERR_INTRO_Q0_0_67_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_67_ERR_INTRO_Q0_0_67_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_68_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_68_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_68_BYTE_OFFSET = 13'h04fc;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_68_ERR_INTRO_Q0_0_68_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_68_ERR_INTRO_Q0_0_68_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_68_ERR_INTRO_Q0_0_68_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_69_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_69_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_69_BYTE_OFFSET = 13'h0500;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_69_ERR_INTRO_Q0_0_69_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_69_ERR_INTRO_Q0_0_69_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_69_ERR_INTRO_Q0_0_69_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_70_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_70_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_70_BYTE_OFFSET = 13'h0504;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_70_ERR_INTRO_Q0_0_70_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_70_ERR_INTRO_Q0_0_70_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_70_ERR_INTRO_Q0_0_70_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_71_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_71_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_71_BYTE_OFFSET = 13'h0508;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_71_ERR_INTRO_Q0_0_71_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_71_ERR_INTRO_Q0_0_71_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_71_ERR_INTRO_Q0_0_71_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_72_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_72_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_72_BYTE_OFFSET = 13'h050c;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_72_ERR_INTRO_Q0_0_72_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_72_ERR_INTRO_Q0_0_72_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_72_ERR_INTRO_Q0_0_72_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_73_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_73_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_73_BYTE_OFFSET = 13'h0510;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_73_ERR_INTRO_Q0_0_73_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_73_ERR_INTRO_Q0_0_73_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_73_ERR_INTRO_Q0_0_73_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_74_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_74_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_74_BYTE_OFFSET = 13'h0514;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_74_ERR_INTRO_Q0_0_74_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_74_ERR_INTRO_Q0_0_74_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_74_ERR_INTRO_Q0_0_74_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_75_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_75_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_75_BYTE_OFFSET = 13'h0518;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_75_ERR_INTRO_Q0_0_75_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_75_ERR_INTRO_Q0_0_75_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_75_ERR_INTRO_Q0_0_75_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_76_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_76_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_76_BYTE_OFFSET = 13'h051c;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_76_ERR_INTRO_Q0_0_76_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_76_ERR_INTRO_Q0_0_76_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_76_ERR_INTRO_Q0_0_76_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_77_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_77_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_77_BYTE_OFFSET = 13'h0520;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_77_ERR_INTRO_Q0_0_77_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_77_ERR_INTRO_Q0_0_77_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_77_ERR_INTRO_Q0_0_77_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_78_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_78_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_78_BYTE_OFFSET = 13'h0524;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_78_ERR_INTRO_Q0_0_78_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_78_ERR_INTRO_Q0_0_78_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_78_ERR_INTRO_Q0_0_78_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_79_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_79_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_79_BYTE_OFFSET = 13'h0528;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_79_ERR_INTRO_Q0_0_79_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_79_ERR_INTRO_Q0_0_79_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_79_ERR_INTRO_Q0_0_79_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_80_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_80_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_80_BYTE_OFFSET = 13'h052c;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_80_ERR_INTRO_Q0_0_80_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_80_ERR_INTRO_Q0_0_80_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_80_ERR_INTRO_Q0_0_80_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_81_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_81_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_81_BYTE_OFFSET = 13'h0530;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_81_ERR_INTRO_Q0_0_81_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_81_ERR_INTRO_Q0_0_81_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_81_ERR_INTRO_Q0_0_81_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_82_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_82_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_82_BYTE_OFFSET = 13'h0534;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_82_ERR_INTRO_Q0_0_82_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_82_ERR_INTRO_Q0_0_82_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_82_ERR_INTRO_Q0_0_82_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_83_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_83_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_83_BYTE_OFFSET = 13'h0538;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_83_ERR_INTRO_Q0_0_83_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_83_ERR_INTRO_Q0_0_83_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_83_ERR_INTRO_Q0_0_83_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_84_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_84_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_84_BYTE_OFFSET = 13'h053c;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_84_ERR_INTRO_Q0_0_84_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_84_ERR_INTRO_Q0_0_84_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_84_ERR_INTRO_Q0_0_84_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_85_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_85_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_85_BYTE_OFFSET = 13'h0540;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_85_ERR_INTRO_Q0_0_85_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_85_ERR_INTRO_Q0_0_85_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_85_ERR_INTRO_Q0_0_85_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_86_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_86_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_86_BYTE_OFFSET = 13'h0544;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_86_ERR_INTRO_Q0_0_86_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_86_ERR_INTRO_Q0_0_86_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_86_ERR_INTRO_Q0_0_86_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_87_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_87_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_87_BYTE_OFFSET = 13'h0548;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_87_ERR_INTRO_Q0_0_87_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_87_ERR_INTRO_Q0_0_87_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_87_ERR_INTRO_Q0_0_87_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_88_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_88_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_88_BYTE_OFFSET = 13'h054c;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_88_ERR_INTRO_Q0_0_88_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_88_ERR_INTRO_Q0_0_88_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_88_ERR_INTRO_Q0_0_88_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_89_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_89_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_89_BYTE_OFFSET = 13'h0550;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_89_ERR_INTRO_Q0_0_89_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_89_ERR_INTRO_Q0_0_89_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_89_ERR_INTRO_Q0_0_89_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_90_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_90_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_90_BYTE_OFFSET = 13'h0554;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_90_ERR_INTRO_Q0_0_90_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_90_ERR_INTRO_Q0_0_90_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_90_ERR_INTRO_Q0_0_90_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_91_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_91_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_91_BYTE_OFFSET = 13'h0558;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_91_ERR_INTRO_Q0_0_91_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_91_ERR_INTRO_Q0_0_91_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_91_ERR_INTRO_Q0_0_91_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_92_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_92_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_92_BYTE_OFFSET = 13'h055c;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_92_ERR_INTRO_Q0_0_92_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_92_ERR_INTRO_Q0_0_92_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_92_ERR_INTRO_Q0_0_92_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_93_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_93_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_93_BYTE_OFFSET = 13'h0560;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_93_ERR_INTRO_Q0_0_93_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_93_ERR_INTRO_Q0_0_93_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_93_ERR_INTRO_Q0_0_93_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_94_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_94_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_94_BYTE_OFFSET = 13'h0564;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_94_ERR_INTRO_Q0_0_94_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_94_ERR_INTRO_Q0_0_94_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_94_ERR_INTRO_Q0_0_94_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_95_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_95_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_95_BYTE_OFFSET = 13'h0568;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_95_ERR_INTRO_Q0_0_95_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_95_ERR_INTRO_Q0_0_95_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_95_ERR_INTRO_Q0_0_95_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_96_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_96_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_96_BYTE_OFFSET = 13'h056c;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_96_ERR_INTRO_Q0_0_96_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_96_ERR_INTRO_Q0_0_96_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_96_ERR_INTRO_Q0_0_96_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_97_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_97_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_97_BYTE_OFFSET = 13'h0570;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_97_ERR_INTRO_Q0_0_97_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_97_ERR_INTRO_Q0_0_97_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_97_ERR_INTRO_Q0_0_97_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_98_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_98_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_98_BYTE_OFFSET = 13'h0574;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_98_ERR_INTRO_Q0_0_98_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_98_ERR_INTRO_Q0_0_98_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_98_ERR_INTRO_Q0_0_98_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_99_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_99_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_99_BYTE_OFFSET = 13'h0578;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_99_ERR_INTRO_Q0_0_99_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_99_ERR_INTRO_Q0_0_99_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_99_ERR_INTRO_Q0_0_99_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_100_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_100_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_100_BYTE_OFFSET = 13'h057c;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_100_ERR_INTRO_Q0_0_100_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_100_ERR_INTRO_Q0_0_100_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_100_ERR_INTRO_Q0_0_100_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_101_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_101_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_101_BYTE_OFFSET = 13'h0580;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_101_ERR_INTRO_Q0_0_101_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_101_ERR_INTRO_Q0_0_101_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_101_ERR_INTRO_Q0_0_101_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_102_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_102_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_102_BYTE_OFFSET = 13'h0584;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_102_ERR_INTRO_Q0_0_102_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_102_ERR_INTRO_Q0_0_102_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_102_ERR_INTRO_Q0_0_102_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_103_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_103_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_103_BYTE_OFFSET = 13'h0588;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_103_ERR_INTRO_Q0_0_103_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_103_ERR_INTRO_Q0_0_103_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_103_ERR_INTRO_Q0_0_103_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_104_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_104_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_104_BYTE_OFFSET = 13'h058c;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_104_ERR_INTRO_Q0_0_104_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_104_ERR_INTRO_Q0_0_104_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_104_ERR_INTRO_Q0_0_104_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_105_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_105_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_105_BYTE_OFFSET = 13'h0590;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_105_ERR_INTRO_Q0_0_105_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_105_ERR_INTRO_Q0_0_105_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_105_ERR_INTRO_Q0_0_105_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_106_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_106_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_106_BYTE_OFFSET = 13'h0594;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_106_ERR_INTRO_Q0_0_106_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_106_ERR_INTRO_Q0_0_106_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_106_ERR_INTRO_Q0_0_106_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_107_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_107_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_107_BYTE_OFFSET = 13'h0598;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_107_ERR_INTRO_Q0_0_107_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_107_ERR_INTRO_Q0_0_107_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_107_ERR_INTRO_Q0_0_107_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_108_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_108_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_108_BYTE_OFFSET = 13'h059c;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_108_ERR_INTRO_Q0_0_108_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_108_ERR_INTRO_Q0_0_108_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_108_ERR_INTRO_Q0_0_108_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_109_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_109_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_109_BYTE_OFFSET = 13'h05a0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_109_ERR_INTRO_Q0_0_109_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_109_ERR_INTRO_Q0_0_109_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_109_ERR_INTRO_Q0_0_109_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_110_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_110_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_110_BYTE_OFFSET = 13'h05a4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_110_ERR_INTRO_Q0_0_110_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_110_ERR_INTRO_Q0_0_110_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_110_ERR_INTRO_Q0_0_110_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_111_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_111_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_111_BYTE_OFFSET = 13'h05a8;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_111_ERR_INTRO_Q0_0_111_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_111_ERR_INTRO_Q0_0_111_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_111_ERR_INTRO_Q0_0_111_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_112_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_112_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_112_BYTE_OFFSET = 13'h05ac;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_112_ERR_INTRO_Q0_0_112_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_112_ERR_INTRO_Q0_0_112_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_112_ERR_INTRO_Q0_0_112_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_113_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_113_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_113_BYTE_OFFSET = 13'h05b0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_113_ERR_INTRO_Q0_0_113_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_113_ERR_INTRO_Q0_0_113_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_113_ERR_INTRO_Q0_0_113_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_114_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_114_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_114_BYTE_OFFSET = 13'h05b4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_114_ERR_INTRO_Q0_0_114_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_114_ERR_INTRO_Q0_0_114_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_114_ERR_INTRO_Q0_0_114_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_115_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_115_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_115_BYTE_OFFSET = 13'h05b8;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_115_ERR_INTRO_Q0_0_115_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_115_ERR_INTRO_Q0_0_115_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_115_ERR_INTRO_Q0_0_115_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_116_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_116_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_116_BYTE_OFFSET = 13'h05bc;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_116_ERR_INTRO_Q0_0_116_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_116_ERR_INTRO_Q0_0_116_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_116_ERR_INTRO_Q0_0_116_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_117_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_117_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_117_BYTE_OFFSET = 13'h05c0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_117_ERR_INTRO_Q0_0_117_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_117_ERR_INTRO_Q0_0_117_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_117_ERR_INTRO_Q0_0_117_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_118_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_118_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_118_BYTE_OFFSET = 13'h05c4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_118_ERR_INTRO_Q0_0_118_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_118_ERR_INTRO_Q0_0_118_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_118_ERR_INTRO_Q0_0_118_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_119_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_119_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_119_BYTE_OFFSET = 13'h05c8;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_119_ERR_INTRO_Q0_0_119_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_119_ERR_INTRO_Q0_0_119_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_119_ERR_INTRO_Q0_0_119_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_120_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_120_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_120_BYTE_OFFSET = 13'h05cc;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_120_ERR_INTRO_Q0_0_120_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_120_ERR_INTRO_Q0_0_120_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_120_ERR_INTRO_Q0_0_120_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_121_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_121_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_121_BYTE_OFFSET = 13'h05d0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_121_ERR_INTRO_Q0_0_121_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_121_ERR_INTRO_Q0_0_121_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_121_ERR_INTRO_Q0_0_121_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_122_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_122_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_122_BYTE_OFFSET = 13'h05d4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_122_ERR_INTRO_Q0_0_122_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_122_ERR_INTRO_Q0_0_122_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_122_ERR_INTRO_Q0_0_122_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_123_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_123_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_123_BYTE_OFFSET = 13'h05d8;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_123_ERR_INTRO_Q0_0_123_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_123_ERR_INTRO_Q0_0_123_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_123_ERR_INTRO_Q0_0_123_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_124_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_124_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_124_BYTE_OFFSET = 13'h05dc;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_124_ERR_INTRO_Q0_0_124_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_124_ERR_INTRO_Q0_0_124_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_124_ERR_INTRO_Q0_0_124_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_125_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_125_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_125_BYTE_OFFSET = 13'h05e0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_125_ERR_INTRO_Q0_0_125_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_125_ERR_INTRO_Q0_0_125_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_125_ERR_INTRO_Q0_0_125_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_126_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_126_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_126_BYTE_OFFSET = 13'h05e4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_126_ERR_INTRO_Q0_0_126_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_126_ERR_INTRO_Q0_0_126_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_126_ERR_INTRO_Q0_0_126_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_127_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_127_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_127_BYTE_OFFSET = 13'h05e8;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_127_ERR_INTRO_Q0_0_127_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_127_ERR_INTRO_Q0_0_127_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_127_ERR_INTRO_Q0_0_127_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_128_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_128_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_128_BYTE_OFFSET = 13'h05ec;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_128_ERR_INTRO_Q0_0_128_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_128_ERR_INTRO_Q0_0_128_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_128_ERR_INTRO_Q0_0_128_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_129_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_129_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_129_BYTE_OFFSET = 13'h05f0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_129_ERR_INTRO_Q0_0_129_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_129_ERR_INTRO_Q0_0_129_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_129_ERR_INTRO_Q0_0_129_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_130_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_130_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_130_BYTE_OFFSET = 13'h05f4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_130_ERR_INTRO_Q0_0_130_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_130_ERR_INTRO_Q0_0_130_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_130_ERR_INTRO_Q0_0_130_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_131_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_131_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_131_BYTE_OFFSET = 13'h05f8;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_131_ERR_INTRO_Q0_0_131_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_131_ERR_INTRO_Q0_0_131_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_131_ERR_INTRO_Q0_0_131_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_132_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_132_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_132_BYTE_OFFSET = 13'h05fc;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_132_ERR_INTRO_Q0_0_132_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_132_ERR_INTRO_Q0_0_132_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_132_ERR_INTRO_Q0_0_132_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_133_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_133_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_133_BYTE_OFFSET = 13'h0600;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_133_ERR_INTRO_Q0_0_133_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_133_ERR_INTRO_Q0_0_133_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_133_ERR_INTRO_Q0_0_133_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_134_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_134_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_134_BYTE_OFFSET = 13'h0604;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_134_ERR_INTRO_Q0_0_134_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_134_ERR_INTRO_Q0_0_134_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_134_ERR_INTRO_Q0_0_134_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_135_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_135_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_135_BYTE_OFFSET = 13'h0608;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_135_ERR_INTRO_Q0_0_135_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_135_ERR_INTRO_Q0_0_135_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_135_ERR_INTRO_Q0_0_135_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_136_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_136_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_136_BYTE_OFFSET = 13'h060c;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_136_ERR_INTRO_Q0_0_136_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_136_ERR_INTRO_Q0_0_136_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_136_ERR_INTRO_Q0_0_136_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_137_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_137_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_137_BYTE_OFFSET = 13'h0610;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_137_ERR_INTRO_Q0_0_137_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_137_ERR_INTRO_Q0_0_137_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_137_ERR_INTRO_Q0_0_137_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_138_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_138_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_138_BYTE_OFFSET = 13'h0614;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_138_ERR_INTRO_Q0_0_138_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_138_ERR_INTRO_Q0_0_138_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_138_ERR_INTRO_Q0_0_138_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_139_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_139_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_139_BYTE_OFFSET = 13'h0618;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_139_ERR_INTRO_Q0_0_139_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_139_ERR_INTRO_Q0_0_139_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_139_ERR_INTRO_Q0_0_139_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_140_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_140_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_140_BYTE_OFFSET = 13'h061c;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_140_ERR_INTRO_Q0_0_140_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_140_ERR_INTRO_Q0_0_140_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_140_ERR_INTRO_Q0_0_140_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_141_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_141_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_141_BYTE_OFFSET = 13'h0620;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_141_ERR_INTRO_Q0_0_141_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_141_ERR_INTRO_Q0_0_141_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_141_ERR_INTRO_Q0_0_141_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_142_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_142_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_142_BYTE_OFFSET = 13'h0624;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_142_ERR_INTRO_Q0_0_142_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_142_ERR_INTRO_Q0_0_142_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_142_ERR_INTRO_Q0_0_142_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_143_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_143_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_143_BYTE_OFFSET = 13'h0628;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_143_ERR_INTRO_Q0_0_143_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_143_ERR_INTRO_Q0_0_143_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_143_ERR_INTRO_Q0_0_143_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_144_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_144_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_144_BYTE_OFFSET = 13'h062c;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_144_ERR_INTRO_Q0_0_144_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_144_ERR_INTRO_Q0_0_144_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_144_ERR_INTRO_Q0_0_144_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_145_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_145_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_145_BYTE_OFFSET = 13'h0630;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_145_ERR_INTRO_Q0_0_145_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_145_ERR_INTRO_Q0_0_145_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_145_ERR_INTRO_Q0_0_145_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_146_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_146_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_146_BYTE_OFFSET = 13'h0634;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_146_ERR_INTRO_Q0_0_146_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_146_ERR_INTRO_Q0_0_146_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_146_ERR_INTRO_Q0_0_146_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_147_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_147_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_147_BYTE_OFFSET = 13'h0638;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_147_ERR_INTRO_Q0_0_147_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_147_ERR_INTRO_Q0_0_147_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_147_ERR_INTRO_Q0_0_147_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_148_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_148_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_148_BYTE_OFFSET = 13'h063c;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_148_ERR_INTRO_Q0_0_148_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_148_ERR_INTRO_Q0_0_148_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_148_ERR_INTRO_Q0_0_148_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_149_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_149_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_149_BYTE_OFFSET = 13'h0640;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_149_ERR_INTRO_Q0_0_149_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_149_ERR_INTRO_Q0_0_149_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_149_ERR_INTRO_Q0_0_149_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_150_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_150_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_150_BYTE_OFFSET = 13'h0644;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_150_ERR_INTRO_Q0_0_150_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_150_ERR_INTRO_Q0_0_150_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_150_ERR_INTRO_Q0_0_150_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_151_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_151_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_151_BYTE_OFFSET = 13'h0648;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_151_ERR_INTRO_Q0_0_151_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_151_ERR_INTRO_Q0_0_151_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_151_ERR_INTRO_Q0_0_151_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_152_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_152_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_152_BYTE_OFFSET = 13'h064c;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_152_ERR_INTRO_Q0_0_152_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_152_ERR_INTRO_Q0_0_152_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_152_ERR_INTRO_Q0_0_152_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_153_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_153_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_153_BYTE_OFFSET = 13'h0650;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_153_ERR_INTRO_Q0_0_153_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_153_ERR_INTRO_Q0_0_153_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_153_ERR_INTRO_Q0_0_153_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_154_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_154_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_154_BYTE_OFFSET = 13'h0654;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_154_ERR_INTRO_Q0_0_154_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_154_ERR_INTRO_Q0_0_154_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_154_ERR_INTRO_Q0_0_154_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_155_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_155_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_155_BYTE_OFFSET = 13'h0658;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_155_ERR_INTRO_Q0_0_155_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_155_ERR_INTRO_Q0_0_155_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_155_ERR_INTRO_Q0_0_155_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_156_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_156_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_156_BYTE_OFFSET = 13'h065c;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_156_ERR_INTRO_Q0_0_156_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_156_ERR_INTRO_Q0_0_156_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_156_ERR_INTRO_Q0_0_156_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_157_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_157_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_157_BYTE_OFFSET = 13'h0660;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_157_ERR_INTRO_Q0_0_157_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_157_ERR_INTRO_Q0_0_157_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_157_ERR_INTRO_Q0_0_157_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_158_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_158_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_158_BYTE_OFFSET = 13'h0664;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_158_ERR_INTRO_Q0_0_158_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_158_ERR_INTRO_Q0_0_158_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_158_ERR_INTRO_Q0_0_158_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_159_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_159_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_159_BYTE_OFFSET = 13'h0668;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_159_ERR_INTRO_Q0_0_159_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_159_ERR_INTRO_Q0_0_159_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_159_ERR_INTRO_Q0_0_159_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_160_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_160_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_160_BYTE_OFFSET = 13'h066c;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_160_ERR_INTRO_Q0_0_160_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_160_ERR_INTRO_Q0_0_160_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_160_ERR_INTRO_Q0_0_160_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_161_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_161_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_161_BYTE_OFFSET = 13'h0670;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_161_ERR_INTRO_Q0_0_161_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_161_ERR_INTRO_Q0_0_161_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_161_ERR_INTRO_Q0_0_161_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_162_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_162_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_162_BYTE_OFFSET = 13'h0674;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_162_ERR_INTRO_Q0_0_162_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_162_ERR_INTRO_Q0_0_162_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_162_ERR_INTRO_Q0_0_162_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_163_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_163_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_163_BYTE_OFFSET = 13'h0678;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_163_ERR_INTRO_Q0_0_163_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_163_ERR_INTRO_Q0_0_163_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_163_ERR_INTRO_Q0_0_163_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_164_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_164_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_164_BYTE_OFFSET = 13'h067c;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_164_ERR_INTRO_Q0_0_164_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_164_ERR_INTRO_Q0_0_164_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_164_ERR_INTRO_Q0_0_164_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_165_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_165_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_165_BYTE_OFFSET = 13'h0680;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_165_ERR_INTRO_Q0_0_165_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_165_ERR_INTRO_Q0_0_165_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_165_ERR_INTRO_Q0_0_165_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_166_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_166_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_166_BYTE_OFFSET = 13'h0684;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_166_ERR_INTRO_Q0_0_166_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_166_ERR_INTRO_Q0_0_166_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_166_ERR_INTRO_Q0_0_166_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_167_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_167_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_167_BYTE_OFFSET = 13'h0688;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_167_ERR_INTRO_Q0_0_167_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_167_ERR_INTRO_Q0_0_167_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_167_ERR_INTRO_Q0_0_167_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_168_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_168_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_168_BYTE_OFFSET = 13'h068c;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_168_ERR_INTRO_Q0_0_168_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_168_ERR_INTRO_Q0_0_168_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_168_ERR_INTRO_Q0_0_168_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_169_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_169_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_169_BYTE_OFFSET = 13'h0690;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_169_ERR_INTRO_Q0_0_169_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_169_ERR_INTRO_Q0_0_169_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_169_ERR_INTRO_Q0_0_169_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_170_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_170_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_170_BYTE_OFFSET = 13'h0694;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_170_ERR_INTRO_Q0_0_170_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_170_ERR_INTRO_Q0_0_170_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_170_ERR_INTRO_Q0_0_170_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_171_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_171_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_171_BYTE_OFFSET = 13'h0698;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_171_ERR_INTRO_Q0_0_171_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_171_ERR_INTRO_Q0_0_171_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_171_ERR_INTRO_Q0_0_171_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_172_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_172_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_172_BYTE_OFFSET = 13'h069c;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_172_ERR_INTRO_Q0_0_172_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_172_ERR_INTRO_Q0_0_172_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_172_ERR_INTRO_Q0_0_172_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_173_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_173_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_173_BYTE_OFFSET = 13'h06a0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_173_ERR_INTRO_Q0_0_173_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_173_ERR_INTRO_Q0_0_173_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_173_ERR_INTRO_Q0_0_173_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_174_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_174_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_174_BYTE_OFFSET = 13'h06a4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_174_ERR_INTRO_Q0_0_174_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_174_ERR_INTRO_Q0_0_174_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_174_ERR_INTRO_Q0_0_174_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_175_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_175_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_175_BYTE_OFFSET = 13'h06a8;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_175_ERR_INTRO_Q0_0_175_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_175_ERR_INTRO_Q0_0_175_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_175_ERR_INTRO_Q0_0_175_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_176_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_176_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_176_BYTE_OFFSET = 13'h06ac;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_176_ERR_INTRO_Q0_0_176_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_176_ERR_INTRO_Q0_0_176_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_176_ERR_INTRO_Q0_0_176_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_177_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_177_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_177_BYTE_OFFSET = 13'h06b0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_177_ERR_INTRO_Q0_0_177_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_177_ERR_INTRO_Q0_0_177_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_177_ERR_INTRO_Q0_0_177_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_178_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_178_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_178_BYTE_OFFSET = 13'h06b4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_178_ERR_INTRO_Q0_0_178_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_178_ERR_INTRO_Q0_0_178_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_178_ERR_INTRO_Q0_0_178_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_179_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_179_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_179_BYTE_OFFSET = 13'h06b8;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_179_ERR_INTRO_Q0_0_179_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_179_ERR_INTRO_Q0_0_179_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_179_ERR_INTRO_Q0_0_179_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_180_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_180_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_180_BYTE_OFFSET = 13'h06bc;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_180_ERR_INTRO_Q0_0_180_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_180_ERR_INTRO_Q0_0_180_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_180_ERR_INTRO_Q0_0_180_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_181_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_181_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_181_BYTE_OFFSET = 13'h06c0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_181_ERR_INTRO_Q0_0_181_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_181_ERR_INTRO_Q0_0_181_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_181_ERR_INTRO_Q0_0_181_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_182_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_182_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_182_BYTE_OFFSET = 13'h06c4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_182_ERR_INTRO_Q0_0_182_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_182_ERR_INTRO_Q0_0_182_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_182_ERR_INTRO_Q0_0_182_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_183_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_183_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_183_BYTE_OFFSET = 13'h06c8;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_183_ERR_INTRO_Q0_0_183_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_183_ERR_INTRO_Q0_0_183_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_183_ERR_INTRO_Q0_0_183_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_184_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_184_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_184_BYTE_OFFSET = 13'h06cc;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_184_ERR_INTRO_Q0_0_184_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_184_ERR_INTRO_Q0_0_184_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_184_ERR_INTRO_Q0_0_184_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_185_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_185_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_185_BYTE_OFFSET = 13'h06d0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_185_ERR_INTRO_Q0_0_185_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_185_ERR_INTRO_Q0_0_185_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_185_ERR_INTRO_Q0_0_185_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_186_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_186_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_186_BYTE_OFFSET = 13'h06d4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_186_ERR_INTRO_Q0_0_186_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_186_ERR_INTRO_Q0_0_186_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_186_ERR_INTRO_Q0_0_186_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_187_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_187_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_187_BYTE_OFFSET = 13'h06d8;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_187_ERR_INTRO_Q0_0_187_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_187_ERR_INTRO_Q0_0_187_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_187_ERR_INTRO_Q0_0_187_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_188_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_188_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_188_BYTE_OFFSET = 13'h06dc;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_188_ERR_INTRO_Q0_0_188_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_188_ERR_INTRO_Q0_0_188_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_188_ERR_INTRO_Q0_0_188_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_189_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_189_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_189_BYTE_OFFSET = 13'h06e0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_189_ERR_INTRO_Q0_0_189_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_189_ERR_INTRO_Q0_0_189_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_189_ERR_INTRO_Q0_0_189_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_190_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_190_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_190_BYTE_OFFSET = 13'h06e4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_190_ERR_INTRO_Q0_0_190_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_190_ERR_INTRO_Q0_0_190_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_190_ERR_INTRO_Q0_0_190_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_191_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_191_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_191_BYTE_OFFSET = 13'h06e8;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_191_ERR_INTRO_Q0_0_191_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_191_ERR_INTRO_Q0_0_191_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_191_ERR_INTRO_Q0_0_191_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_192_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_192_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_192_BYTE_OFFSET = 13'h06ec;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_192_ERR_INTRO_Q0_0_192_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_192_ERR_INTRO_Q0_0_192_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_192_ERR_INTRO_Q0_0_192_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_193_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_193_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_193_BYTE_OFFSET = 13'h06f0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_193_ERR_INTRO_Q0_0_193_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_193_ERR_INTRO_Q0_0_193_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_193_ERR_INTRO_Q0_0_193_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_194_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_194_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_194_BYTE_OFFSET = 13'h06f4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_194_ERR_INTRO_Q0_0_194_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_194_ERR_INTRO_Q0_0_194_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_194_ERR_INTRO_Q0_0_194_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_195_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_195_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_195_BYTE_OFFSET = 13'h06f8;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_195_ERR_INTRO_Q0_0_195_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_195_ERR_INTRO_Q0_0_195_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_195_ERR_INTRO_Q0_0_195_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_196_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_196_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_196_BYTE_OFFSET = 13'h06fc;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_196_ERR_INTRO_Q0_0_196_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_196_ERR_INTRO_Q0_0_196_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_196_ERR_INTRO_Q0_0_196_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_197_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_197_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_197_BYTE_OFFSET = 13'h0700;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_197_ERR_INTRO_Q0_0_197_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_197_ERR_INTRO_Q0_0_197_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_197_ERR_INTRO_Q0_0_197_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_198_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_198_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_198_BYTE_OFFSET = 13'h0704;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_198_ERR_INTRO_Q0_0_198_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_198_ERR_INTRO_Q0_0_198_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_198_ERR_INTRO_Q0_0_198_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_199_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_199_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_199_BYTE_OFFSET = 13'h0708;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_199_ERR_INTRO_Q0_0_199_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_199_ERR_INTRO_Q0_0_199_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_199_ERR_INTRO_Q0_0_199_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_200_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_200_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_200_BYTE_OFFSET = 13'h070c;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_200_ERR_INTRO_Q0_0_200_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_200_ERR_INTRO_Q0_0_200_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_200_ERR_INTRO_Q0_0_200_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_201_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_201_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_201_BYTE_OFFSET = 13'h0710;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_201_ERR_INTRO_Q0_0_201_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_201_ERR_INTRO_Q0_0_201_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_201_ERR_INTRO_Q0_0_201_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_202_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_202_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_202_BYTE_OFFSET = 13'h0714;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_202_ERR_INTRO_Q0_0_202_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_202_ERR_INTRO_Q0_0_202_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_202_ERR_INTRO_Q0_0_202_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_203_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_203_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_203_BYTE_OFFSET = 13'h0718;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_203_ERR_INTRO_Q0_0_203_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_203_ERR_INTRO_Q0_0_203_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_203_ERR_INTRO_Q0_0_203_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_204_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_204_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_204_BYTE_OFFSET = 13'h071c;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_204_ERR_INTRO_Q0_0_204_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_204_ERR_INTRO_Q0_0_204_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_204_ERR_INTRO_Q0_0_204_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_205_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_205_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_205_BYTE_OFFSET = 13'h0720;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_205_ERR_INTRO_Q0_0_205_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_205_ERR_INTRO_Q0_0_205_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_205_ERR_INTRO_Q0_0_205_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_206_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_206_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_206_BYTE_OFFSET = 13'h0724;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_206_ERR_INTRO_Q0_0_206_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_206_ERR_INTRO_Q0_0_206_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_206_ERR_INTRO_Q0_0_206_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_207_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_207_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_0_INTRO_207_BYTE_OFFSET = 13'h0728;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_207_ERR_INTRO_Q0_0_207_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_0_INTRO_207_ERR_INTRO_Q0_0_207_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_0_INTRO_207_ERR_INTRO_Q0_0_207_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_0_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_0_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_0_BYTE_OFFSET = 13'h072c;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_0_ERR_INTRO_Q0_1_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_0_ERR_INTRO_Q0_1_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_0_ERR_INTRO_Q0_1_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_1_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_1_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_1_BYTE_OFFSET = 13'h0730;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_1_ERR_INTRO_Q0_1_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_1_ERR_INTRO_Q0_1_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_1_ERR_INTRO_Q0_1_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_2_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_2_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_2_BYTE_OFFSET = 13'h0734;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_2_ERR_INTRO_Q0_1_2_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_2_ERR_INTRO_Q0_1_2_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_2_ERR_INTRO_Q0_1_2_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_3_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_3_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_3_BYTE_OFFSET = 13'h0738;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_3_ERR_INTRO_Q0_1_3_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_3_ERR_INTRO_Q0_1_3_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_3_ERR_INTRO_Q0_1_3_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_4_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_4_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_4_BYTE_OFFSET = 13'h073c;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_4_ERR_INTRO_Q0_1_4_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_4_ERR_INTRO_Q0_1_4_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_4_ERR_INTRO_Q0_1_4_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_5_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_5_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_5_BYTE_OFFSET = 13'h0740;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_5_ERR_INTRO_Q0_1_5_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_5_ERR_INTRO_Q0_1_5_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_5_ERR_INTRO_Q0_1_5_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_6_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_6_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_6_BYTE_OFFSET = 13'h0744;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_6_ERR_INTRO_Q0_1_6_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_6_ERR_INTRO_Q0_1_6_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_6_ERR_INTRO_Q0_1_6_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_7_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_7_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_7_BYTE_OFFSET = 13'h0748;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_7_ERR_INTRO_Q0_1_7_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_7_ERR_INTRO_Q0_1_7_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_7_ERR_INTRO_Q0_1_7_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_8_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_8_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_8_BYTE_OFFSET = 13'h074c;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_8_ERR_INTRO_Q0_1_8_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_8_ERR_INTRO_Q0_1_8_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_8_ERR_INTRO_Q0_1_8_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_9_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_9_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_9_BYTE_OFFSET = 13'h0750;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_9_ERR_INTRO_Q0_1_9_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_9_ERR_INTRO_Q0_1_9_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_9_ERR_INTRO_Q0_1_9_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_10_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_10_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_10_BYTE_OFFSET = 13'h0754;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_10_ERR_INTRO_Q0_1_10_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_10_ERR_INTRO_Q0_1_10_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_10_ERR_INTRO_Q0_1_10_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_11_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_11_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_11_BYTE_OFFSET = 13'h0758;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_11_ERR_INTRO_Q0_1_11_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_11_ERR_INTRO_Q0_1_11_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_11_ERR_INTRO_Q0_1_11_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_12_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_12_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_12_BYTE_OFFSET = 13'h075c;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_12_ERR_INTRO_Q0_1_12_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_12_ERR_INTRO_Q0_1_12_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_12_ERR_INTRO_Q0_1_12_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_13_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_13_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_13_BYTE_OFFSET = 13'h0760;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_13_ERR_INTRO_Q0_1_13_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_13_ERR_INTRO_Q0_1_13_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_13_ERR_INTRO_Q0_1_13_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_14_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_14_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_14_BYTE_OFFSET = 13'h0764;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_14_ERR_INTRO_Q0_1_14_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_14_ERR_INTRO_Q0_1_14_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_14_ERR_INTRO_Q0_1_14_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_15_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_15_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_15_BYTE_OFFSET = 13'h0768;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_15_ERR_INTRO_Q0_1_15_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_15_ERR_INTRO_Q0_1_15_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_15_ERR_INTRO_Q0_1_15_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_16_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_16_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_16_BYTE_OFFSET = 13'h076c;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_16_ERR_INTRO_Q0_1_16_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_16_ERR_INTRO_Q0_1_16_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_16_ERR_INTRO_Q0_1_16_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_17_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_17_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_17_BYTE_OFFSET = 13'h0770;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_17_ERR_INTRO_Q0_1_17_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_17_ERR_INTRO_Q0_1_17_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_17_ERR_INTRO_Q0_1_17_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_18_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_18_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_18_BYTE_OFFSET = 13'h0774;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_18_ERR_INTRO_Q0_1_18_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_18_ERR_INTRO_Q0_1_18_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_18_ERR_INTRO_Q0_1_18_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_19_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_19_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_19_BYTE_OFFSET = 13'h0778;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_19_ERR_INTRO_Q0_1_19_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_19_ERR_INTRO_Q0_1_19_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_19_ERR_INTRO_Q0_1_19_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_20_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_20_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_20_BYTE_OFFSET = 13'h077c;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_20_ERR_INTRO_Q0_1_20_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_20_ERR_INTRO_Q0_1_20_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_20_ERR_INTRO_Q0_1_20_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_21_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_21_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_21_BYTE_OFFSET = 13'h0780;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_21_ERR_INTRO_Q0_1_21_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_21_ERR_INTRO_Q0_1_21_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_21_ERR_INTRO_Q0_1_21_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_22_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_22_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_22_BYTE_OFFSET = 13'h0784;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_22_ERR_INTRO_Q0_1_22_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_22_ERR_INTRO_Q0_1_22_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_22_ERR_INTRO_Q0_1_22_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_23_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_23_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_23_BYTE_OFFSET = 13'h0788;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_23_ERR_INTRO_Q0_1_23_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_23_ERR_INTRO_Q0_1_23_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_23_ERR_INTRO_Q0_1_23_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_24_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_24_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_24_BYTE_OFFSET = 13'h078c;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_24_ERR_INTRO_Q0_1_24_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_24_ERR_INTRO_Q0_1_24_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_24_ERR_INTRO_Q0_1_24_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_25_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_25_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_25_BYTE_OFFSET = 13'h0790;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_25_ERR_INTRO_Q0_1_25_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_25_ERR_INTRO_Q0_1_25_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_25_ERR_INTRO_Q0_1_25_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_26_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_26_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_26_BYTE_OFFSET = 13'h0794;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_26_ERR_INTRO_Q0_1_26_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_26_ERR_INTRO_Q0_1_26_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_26_ERR_INTRO_Q0_1_26_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_27_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_27_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_27_BYTE_OFFSET = 13'h0798;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_27_ERR_INTRO_Q0_1_27_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_27_ERR_INTRO_Q0_1_27_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_27_ERR_INTRO_Q0_1_27_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_28_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_28_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_28_BYTE_OFFSET = 13'h079c;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_28_ERR_INTRO_Q0_1_28_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_28_ERR_INTRO_Q0_1_28_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_28_ERR_INTRO_Q0_1_28_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_29_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_29_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_29_BYTE_OFFSET = 13'h07a0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_29_ERR_INTRO_Q0_1_29_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_29_ERR_INTRO_Q0_1_29_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_29_ERR_INTRO_Q0_1_29_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_30_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_30_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_30_BYTE_OFFSET = 13'h07a4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_30_ERR_INTRO_Q0_1_30_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_30_ERR_INTRO_Q0_1_30_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_30_ERR_INTRO_Q0_1_30_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_31_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_31_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_31_BYTE_OFFSET = 13'h07a8;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_31_ERR_INTRO_Q0_1_31_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_31_ERR_INTRO_Q0_1_31_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_31_ERR_INTRO_Q0_1_31_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_32_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_32_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_32_BYTE_OFFSET = 13'h07ac;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_32_ERR_INTRO_Q0_1_32_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_32_ERR_INTRO_Q0_1_32_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_32_ERR_INTRO_Q0_1_32_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_33_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_33_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_33_BYTE_OFFSET = 13'h07b0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_33_ERR_INTRO_Q0_1_33_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_33_ERR_INTRO_Q0_1_33_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_33_ERR_INTRO_Q0_1_33_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_34_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_34_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_34_BYTE_OFFSET = 13'h07b4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_34_ERR_INTRO_Q0_1_34_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_34_ERR_INTRO_Q0_1_34_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_34_ERR_INTRO_Q0_1_34_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_35_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_35_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_35_BYTE_OFFSET = 13'h07b8;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_35_ERR_INTRO_Q0_1_35_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_35_ERR_INTRO_Q0_1_35_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_35_ERR_INTRO_Q0_1_35_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_36_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_36_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_36_BYTE_OFFSET = 13'h07bc;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_36_ERR_INTRO_Q0_1_36_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_36_ERR_INTRO_Q0_1_36_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_36_ERR_INTRO_Q0_1_36_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_37_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_37_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_37_BYTE_OFFSET = 13'h07c0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_37_ERR_INTRO_Q0_1_37_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_37_ERR_INTRO_Q0_1_37_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_37_ERR_INTRO_Q0_1_37_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_38_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_38_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_38_BYTE_OFFSET = 13'h07c4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_38_ERR_INTRO_Q0_1_38_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_38_ERR_INTRO_Q0_1_38_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_38_ERR_INTRO_Q0_1_38_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_39_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_39_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_39_BYTE_OFFSET = 13'h07c8;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_39_ERR_INTRO_Q0_1_39_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_39_ERR_INTRO_Q0_1_39_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_39_ERR_INTRO_Q0_1_39_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_40_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_40_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_40_BYTE_OFFSET = 13'h07cc;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_40_ERR_INTRO_Q0_1_40_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_40_ERR_INTRO_Q0_1_40_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_40_ERR_INTRO_Q0_1_40_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_41_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_41_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_41_BYTE_OFFSET = 13'h07d0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_41_ERR_INTRO_Q0_1_41_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_41_ERR_INTRO_Q0_1_41_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_41_ERR_INTRO_Q0_1_41_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_42_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_42_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_42_BYTE_OFFSET = 13'h07d4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_42_ERR_INTRO_Q0_1_42_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_42_ERR_INTRO_Q0_1_42_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_42_ERR_INTRO_Q0_1_42_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_43_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_43_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_43_BYTE_OFFSET = 13'h07d8;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_43_ERR_INTRO_Q0_1_43_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_43_ERR_INTRO_Q0_1_43_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_43_ERR_INTRO_Q0_1_43_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_44_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_44_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_44_BYTE_OFFSET = 13'h07dc;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_44_ERR_INTRO_Q0_1_44_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_44_ERR_INTRO_Q0_1_44_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_44_ERR_INTRO_Q0_1_44_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_45_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_45_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_45_BYTE_OFFSET = 13'h07e0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_45_ERR_INTRO_Q0_1_45_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_45_ERR_INTRO_Q0_1_45_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_45_ERR_INTRO_Q0_1_45_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_46_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_46_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_46_BYTE_OFFSET = 13'h07e4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_46_ERR_INTRO_Q0_1_46_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_46_ERR_INTRO_Q0_1_46_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_46_ERR_INTRO_Q0_1_46_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_47_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_47_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_47_BYTE_OFFSET = 13'h07e8;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_47_ERR_INTRO_Q0_1_47_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_47_ERR_INTRO_Q0_1_47_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_47_ERR_INTRO_Q0_1_47_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_48_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_48_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_48_BYTE_OFFSET = 13'h07ec;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_48_ERR_INTRO_Q0_1_48_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_48_ERR_INTRO_Q0_1_48_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_48_ERR_INTRO_Q0_1_48_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_49_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_49_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_49_BYTE_OFFSET = 13'h07f0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_49_ERR_INTRO_Q0_1_49_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_49_ERR_INTRO_Q0_1_49_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_49_ERR_INTRO_Q0_1_49_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_50_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_50_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_50_BYTE_OFFSET = 13'h07f4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_50_ERR_INTRO_Q0_1_50_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_50_ERR_INTRO_Q0_1_50_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_50_ERR_INTRO_Q0_1_50_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_51_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_51_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_51_BYTE_OFFSET = 13'h07f8;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_51_ERR_INTRO_Q0_1_51_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_51_ERR_INTRO_Q0_1_51_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_51_ERR_INTRO_Q0_1_51_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_52_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_52_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_52_BYTE_OFFSET = 13'h07fc;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_52_ERR_INTRO_Q0_1_52_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_52_ERR_INTRO_Q0_1_52_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_52_ERR_INTRO_Q0_1_52_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_53_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_53_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_53_BYTE_OFFSET = 13'h0800;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_53_ERR_INTRO_Q0_1_53_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_53_ERR_INTRO_Q0_1_53_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_53_ERR_INTRO_Q0_1_53_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_54_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_54_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_54_BYTE_OFFSET = 13'h0804;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_54_ERR_INTRO_Q0_1_54_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_54_ERR_INTRO_Q0_1_54_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_54_ERR_INTRO_Q0_1_54_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_55_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_55_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_55_BYTE_OFFSET = 13'h0808;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_55_ERR_INTRO_Q0_1_55_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_55_ERR_INTRO_Q0_1_55_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_55_ERR_INTRO_Q0_1_55_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_56_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_56_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_56_BYTE_OFFSET = 13'h080c;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_56_ERR_INTRO_Q0_1_56_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_56_ERR_INTRO_Q0_1_56_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_56_ERR_INTRO_Q0_1_56_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_57_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_57_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_57_BYTE_OFFSET = 13'h0810;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_57_ERR_INTRO_Q0_1_57_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_57_ERR_INTRO_Q0_1_57_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_57_ERR_INTRO_Q0_1_57_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_58_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_58_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_58_BYTE_OFFSET = 13'h0814;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_58_ERR_INTRO_Q0_1_58_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_58_ERR_INTRO_Q0_1_58_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_58_ERR_INTRO_Q0_1_58_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_59_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_59_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_59_BYTE_OFFSET = 13'h0818;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_59_ERR_INTRO_Q0_1_59_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_59_ERR_INTRO_Q0_1_59_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_59_ERR_INTRO_Q0_1_59_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_60_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_60_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_60_BYTE_OFFSET = 13'h081c;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_60_ERR_INTRO_Q0_1_60_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_60_ERR_INTRO_Q0_1_60_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_60_ERR_INTRO_Q0_1_60_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_61_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_61_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_61_BYTE_OFFSET = 13'h0820;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_61_ERR_INTRO_Q0_1_61_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_61_ERR_INTRO_Q0_1_61_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_61_ERR_INTRO_Q0_1_61_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_62_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_62_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_62_BYTE_OFFSET = 13'h0824;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_62_ERR_INTRO_Q0_1_62_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_62_ERR_INTRO_Q0_1_62_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_62_ERR_INTRO_Q0_1_62_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_63_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_63_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_63_BYTE_OFFSET = 13'h0828;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_63_ERR_INTRO_Q0_1_63_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_63_ERR_INTRO_Q0_1_63_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_63_ERR_INTRO_Q0_1_63_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_64_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_64_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_64_BYTE_OFFSET = 13'h082c;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_64_ERR_INTRO_Q0_1_64_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_64_ERR_INTRO_Q0_1_64_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_64_ERR_INTRO_Q0_1_64_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_65_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_65_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_65_BYTE_OFFSET = 13'h0830;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_65_ERR_INTRO_Q0_1_65_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_65_ERR_INTRO_Q0_1_65_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_65_ERR_INTRO_Q0_1_65_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_66_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_66_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_66_BYTE_OFFSET = 13'h0834;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_66_ERR_INTRO_Q0_1_66_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_66_ERR_INTRO_Q0_1_66_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_66_ERR_INTRO_Q0_1_66_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_67_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_67_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_67_BYTE_OFFSET = 13'h0838;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_67_ERR_INTRO_Q0_1_67_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_67_ERR_INTRO_Q0_1_67_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_67_ERR_INTRO_Q0_1_67_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_68_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_68_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_68_BYTE_OFFSET = 13'h083c;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_68_ERR_INTRO_Q0_1_68_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_68_ERR_INTRO_Q0_1_68_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_68_ERR_INTRO_Q0_1_68_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_69_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_69_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_69_BYTE_OFFSET = 13'h0840;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_69_ERR_INTRO_Q0_1_69_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_69_ERR_INTRO_Q0_1_69_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_69_ERR_INTRO_Q0_1_69_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_70_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_70_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_70_BYTE_OFFSET = 13'h0844;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_70_ERR_INTRO_Q0_1_70_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_70_ERR_INTRO_Q0_1_70_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_70_ERR_INTRO_Q0_1_70_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_71_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_71_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_71_BYTE_OFFSET = 13'h0848;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_71_ERR_INTRO_Q0_1_71_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_71_ERR_INTRO_Q0_1_71_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_71_ERR_INTRO_Q0_1_71_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_72_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_72_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_72_BYTE_OFFSET = 13'h084c;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_72_ERR_INTRO_Q0_1_72_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_72_ERR_INTRO_Q0_1_72_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_72_ERR_INTRO_Q0_1_72_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_73_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_73_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_73_BYTE_OFFSET = 13'h0850;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_73_ERR_INTRO_Q0_1_73_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_73_ERR_INTRO_Q0_1_73_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_73_ERR_INTRO_Q0_1_73_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_74_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_74_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_74_BYTE_OFFSET = 13'h0854;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_74_ERR_INTRO_Q0_1_74_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_74_ERR_INTRO_Q0_1_74_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_74_ERR_INTRO_Q0_1_74_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_75_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_75_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_75_BYTE_OFFSET = 13'h0858;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_75_ERR_INTRO_Q0_1_75_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_75_ERR_INTRO_Q0_1_75_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_75_ERR_INTRO_Q0_1_75_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_76_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_76_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_76_BYTE_OFFSET = 13'h085c;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_76_ERR_INTRO_Q0_1_76_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_76_ERR_INTRO_Q0_1_76_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_76_ERR_INTRO_Q0_1_76_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_77_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_77_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_77_BYTE_OFFSET = 13'h0860;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_77_ERR_INTRO_Q0_1_77_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_77_ERR_INTRO_Q0_1_77_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_77_ERR_INTRO_Q0_1_77_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_78_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_78_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_78_BYTE_OFFSET = 13'h0864;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_78_ERR_INTRO_Q0_1_78_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_78_ERR_INTRO_Q0_1_78_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_78_ERR_INTRO_Q0_1_78_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_79_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_79_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_79_BYTE_OFFSET = 13'h0868;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_79_ERR_INTRO_Q0_1_79_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_79_ERR_INTRO_Q0_1_79_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_79_ERR_INTRO_Q0_1_79_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_80_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_80_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_80_BYTE_OFFSET = 13'h086c;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_80_ERR_INTRO_Q0_1_80_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_80_ERR_INTRO_Q0_1_80_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_80_ERR_INTRO_Q0_1_80_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_81_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_81_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_81_BYTE_OFFSET = 13'h0870;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_81_ERR_INTRO_Q0_1_81_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_81_ERR_INTRO_Q0_1_81_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_81_ERR_INTRO_Q0_1_81_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_82_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_82_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_82_BYTE_OFFSET = 13'h0874;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_82_ERR_INTRO_Q0_1_82_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_82_ERR_INTRO_Q0_1_82_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_82_ERR_INTRO_Q0_1_82_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_83_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_83_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_83_BYTE_OFFSET = 13'h0878;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_83_ERR_INTRO_Q0_1_83_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_83_ERR_INTRO_Q0_1_83_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_83_ERR_INTRO_Q0_1_83_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_84_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_84_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_84_BYTE_OFFSET = 13'h087c;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_84_ERR_INTRO_Q0_1_84_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_84_ERR_INTRO_Q0_1_84_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_84_ERR_INTRO_Q0_1_84_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_85_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_85_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_85_BYTE_OFFSET = 13'h0880;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_85_ERR_INTRO_Q0_1_85_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_85_ERR_INTRO_Q0_1_85_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_85_ERR_INTRO_Q0_1_85_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_86_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_86_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_86_BYTE_OFFSET = 13'h0884;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_86_ERR_INTRO_Q0_1_86_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_86_ERR_INTRO_Q0_1_86_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_86_ERR_INTRO_Q0_1_86_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_87_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_87_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_87_BYTE_OFFSET = 13'h0888;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_87_ERR_INTRO_Q0_1_87_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_87_ERR_INTRO_Q0_1_87_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_87_ERR_INTRO_Q0_1_87_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_88_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_88_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_88_BYTE_OFFSET = 13'h088c;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_88_ERR_INTRO_Q0_1_88_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_88_ERR_INTRO_Q0_1_88_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_88_ERR_INTRO_Q0_1_88_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_89_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_89_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_89_BYTE_OFFSET = 13'h0890;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_89_ERR_INTRO_Q0_1_89_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_89_ERR_INTRO_Q0_1_89_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_89_ERR_INTRO_Q0_1_89_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_90_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_90_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_90_BYTE_OFFSET = 13'h0894;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_90_ERR_INTRO_Q0_1_90_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_90_ERR_INTRO_Q0_1_90_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_90_ERR_INTRO_Q0_1_90_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_91_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_91_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_91_BYTE_OFFSET = 13'h0898;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_91_ERR_INTRO_Q0_1_91_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_91_ERR_INTRO_Q0_1_91_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_91_ERR_INTRO_Q0_1_91_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_92_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_92_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_92_BYTE_OFFSET = 13'h089c;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_92_ERR_INTRO_Q0_1_92_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_92_ERR_INTRO_Q0_1_92_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_92_ERR_INTRO_Q0_1_92_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_93_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_93_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_93_BYTE_OFFSET = 13'h08a0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_93_ERR_INTRO_Q0_1_93_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_93_ERR_INTRO_Q0_1_93_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_93_ERR_INTRO_Q0_1_93_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_94_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_94_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_94_BYTE_OFFSET = 13'h08a4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_94_ERR_INTRO_Q0_1_94_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_94_ERR_INTRO_Q0_1_94_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_94_ERR_INTRO_Q0_1_94_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_95_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_95_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_95_BYTE_OFFSET = 13'h08a8;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_95_ERR_INTRO_Q0_1_95_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_95_ERR_INTRO_Q0_1_95_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_95_ERR_INTRO_Q0_1_95_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_96_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_96_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_96_BYTE_OFFSET = 13'h08ac;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_96_ERR_INTRO_Q0_1_96_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_96_ERR_INTRO_Q0_1_96_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_96_ERR_INTRO_Q0_1_96_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_97_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_97_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_97_BYTE_OFFSET = 13'h08b0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_97_ERR_INTRO_Q0_1_97_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_97_ERR_INTRO_Q0_1_97_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_97_ERR_INTRO_Q0_1_97_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_98_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_98_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_98_BYTE_OFFSET = 13'h08b4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_98_ERR_INTRO_Q0_1_98_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_98_ERR_INTRO_Q0_1_98_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_98_ERR_INTRO_Q0_1_98_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_99_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_99_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_99_BYTE_OFFSET = 13'h08b8;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_99_ERR_INTRO_Q0_1_99_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_99_ERR_INTRO_Q0_1_99_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_99_ERR_INTRO_Q0_1_99_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_100_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_100_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_100_BYTE_OFFSET = 13'h08bc;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_100_ERR_INTRO_Q0_1_100_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_100_ERR_INTRO_Q0_1_100_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_100_ERR_INTRO_Q0_1_100_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_101_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_101_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_101_BYTE_OFFSET = 13'h08c0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_101_ERR_INTRO_Q0_1_101_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_101_ERR_INTRO_Q0_1_101_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_101_ERR_INTRO_Q0_1_101_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_102_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_102_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_102_BYTE_OFFSET = 13'h08c4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_102_ERR_INTRO_Q0_1_102_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_102_ERR_INTRO_Q0_1_102_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_102_ERR_INTRO_Q0_1_102_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_103_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_103_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_103_BYTE_OFFSET = 13'h08c8;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_103_ERR_INTRO_Q0_1_103_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_103_ERR_INTRO_Q0_1_103_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_103_ERR_INTRO_Q0_1_103_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_104_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_104_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_104_BYTE_OFFSET = 13'h08cc;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_104_ERR_INTRO_Q0_1_104_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_104_ERR_INTRO_Q0_1_104_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_104_ERR_INTRO_Q0_1_104_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_105_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_105_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_105_BYTE_OFFSET = 13'h08d0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_105_ERR_INTRO_Q0_1_105_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_105_ERR_INTRO_Q0_1_105_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_105_ERR_INTRO_Q0_1_105_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_106_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_106_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_106_BYTE_OFFSET = 13'h08d4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_106_ERR_INTRO_Q0_1_106_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_106_ERR_INTRO_Q0_1_106_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_106_ERR_INTRO_Q0_1_106_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_107_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_107_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_107_BYTE_OFFSET = 13'h08d8;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_107_ERR_INTRO_Q0_1_107_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_107_ERR_INTRO_Q0_1_107_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_107_ERR_INTRO_Q0_1_107_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_108_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_108_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_108_BYTE_OFFSET = 13'h08dc;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_108_ERR_INTRO_Q0_1_108_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_108_ERR_INTRO_Q0_1_108_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_108_ERR_INTRO_Q0_1_108_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_109_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_109_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_109_BYTE_OFFSET = 13'h08e0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_109_ERR_INTRO_Q0_1_109_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_109_ERR_INTRO_Q0_1_109_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_109_ERR_INTRO_Q0_1_109_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_110_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_110_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_110_BYTE_OFFSET = 13'h08e4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_110_ERR_INTRO_Q0_1_110_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_110_ERR_INTRO_Q0_1_110_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_110_ERR_INTRO_Q0_1_110_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_111_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_111_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_111_BYTE_OFFSET = 13'h08e8;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_111_ERR_INTRO_Q0_1_111_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_111_ERR_INTRO_Q0_1_111_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_111_ERR_INTRO_Q0_1_111_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_112_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_112_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_112_BYTE_OFFSET = 13'h08ec;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_112_ERR_INTRO_Q0_1_112_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_112_ERR_INTRO_Q0_1_112_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_112_ERR_INTRO_Q0_1_112_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_113_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_113_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_113_BYTE_OFFSET = 13'h08f0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_113_ERR_INTRO_Q0_1_113_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_113_ERR_INTRO_Q0_1_113_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_113_ERR_INTRO_Q0_1_113_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_114_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_114_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_114_BYTE_OFFSET = 13'h08f4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_114_ERR_INTRO_Q0_1_114_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_114_ERR_INTRO_Q0_1_114_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_114_ERR_INTRO_Q0_1_114_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_115_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_115_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_115_BYTE_OFFSET = 13'h08f8;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_115_ERR_INTRO_Q0_1_115_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_115_ERR_INTRO_Q0_1_115_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_115_ERR_INTRO_Q0_1_115_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_116_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_116_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_116_BYTE_OFFSET = 13'h08fc;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_116_ERR_INTRO_Q0_1_116_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_116_ERR_INTRO_Q0_1_116_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_116_ERR_INTRO_Q0_1_116_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_117_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_117_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_117_BYTE_OFFSET = 13'h0900;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_117_ERR_INTRO_Q0_1_117_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_117_ERR_INTRO_Q0_1_117_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_117_ERR_INTRO_Q0_1_117_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_118_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_118_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_118_BYTE_OFFSET = 13'h0904;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_118_ERR_INTRO_Q0_1_118_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_118_ERR_INTRO_Q0_1_118_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_118_ERR_INTRO_Q0_1_118_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_119_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_119_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_119_BYTE_OFFSET = 13'h0908;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_119_ERR_INTRO_Q0_1_119_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_119_ERR_INTRO_Q0_1_119_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_119_ERR_INTRO_Q0_1_119_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_120_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_120_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_120_BYTE_OFFSET = 13'h090c;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_120_ERR_INTRO_Q0_1_120_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_120_ERR_INTRO_Q0_1_120_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_120_ERR_INTRO_Q0_1_120_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_121_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_121_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_121_BYTE_OFFSET = 13'h0910;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_121_ERR_INTRO_Q0_1_121_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_121_ERR_INTRO_Q0_1_121_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_121_ERR_INTRO_Q0_1_121_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_122_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_122_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_122_BYTE_OFFSET = 13'h0914;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_122_ERR_INTRO_Q0_1_122_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_122_ERR_INTRO_Q0_1_122_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_122_ERR_INTRO_Q0_1_122_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_123_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_123_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_123_BYTE_OFFSET = 13'h0918;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_123_ERR_INTRO_Q0_1_123_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_123_ERR_INTRO_Q0_1_123_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_123_ERR_INTRO_Q0_1_123_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_124_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_124_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_124_BYTE_OFFSET = 13'h091c;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_124_ERR_INTRO_Q0_1_124_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_124_ERR_INTRO_Q0_1_124_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_124_ERR_INTRO_Q0_1_124_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_125_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_125_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_125_BYTE_OFFSET = 13'h0920;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_125_ERR_INTRO_Q0_1_125_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_125_ERR_INTRO_Q0_1_125_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_125_ERR_INTRO_Q0_1_125_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_126_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_126_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_126_BYTE_OFFSET = 13'h0924;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_126_ERR_INTRO_Q0_1_126_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_126_ERR_INTRO_Q0_1_126_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_126_ERR_INTRO_Q0_1_126_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_127_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_127_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_127_BYTE_OFFSET = 13'h0928;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_127_ERR_INTRO_Q0_1_127_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_127_ERR_INTRO_Q0_1_127_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_127_ERR_INTRO_Q0_1_127_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_128_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_128_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_128_BYTE_OFFSET = 13'h092c;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_128_ERR_INTRO_Q0_1_128_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_128_ERR_INTRO_Q0_1_128_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_128_ERR_INTRO_Q0_1_128_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_129_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_129_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_129_BYTE_OFFSET = 13'h0930;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_129_ERR_INTRO_Q0_1_129_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_129_ERR_INTRO_Q0_1_129_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_129_ERR_INTRO_Q0_1_129_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_130_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_130_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_130_BYTE_OFFSET = 13'h0934;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_130_ERR_INTRO_Q0_1_130_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_130_ERR_INTRO_Q0_1_130_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_130_ERR_INTRO_Q0_1_130_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_131_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_131_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_131_BYTE_OFFSET = 13'h0938;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_131_ERR_INTRO_Q0_1_131_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_131_ERR_INTRO_Q0_1_131_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_131_ERR_INTRO_Q0_1_131_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_132_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_132_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_132_BYTE_OFFSET = 13'h093c;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_132_ERR_INTRO_Q0_1_132_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_132_ERR_INTRO_Q0_1_132_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_132_ERR_INTRO_Q0_1_132_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_133_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_133_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_133_BYTE_OFFSET = 13'h0940;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_133_ERR_INTRO_Q0_1_133_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_133_ERR_INTRO_Q0_1_133_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_133_ERR_INTRO_Q0_1_133_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_134_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_134_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_134_BYTE_OFFSET = 13'h0944;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_134_ERR_INTRO_Q0_1_134_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_134_ERR_INTRO_Q0_1_134_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_134_ERR_INTRO_Q0_1_134_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_135_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_135_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_135_BYTE_OFFSET = 13'h0948;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_135_ERR_INTRO_Q0_1_135_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_135_ERR_INTRO_Q0_1_135_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_135_ERR_INTRO_Q0_1_135_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_136_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_136_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_136_BYTE_OFFSET = 13'h094c;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_136_ERR_INTRO_Q0_1_136_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_136_ERR_INTRO_Q0_1_136_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_136_ERR_INTRO_Q0_1_136_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_137_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_137_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_137_BYTE_OFFSET = 13'h0950;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_137_ERR_INTRO_Q0_1_137_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_137_ERR_INTRO_Q0_1_137_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_137_ERR_INTRO_Q0_1_137_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_138_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_138_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_138_BYTE_OFFSET = 13'h0954;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_138_ERR_INTRO_Q0_1_138_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_138_ERR_INTRO_Q0_1_138_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_138_ERR_INTRO_Q0_1_138_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_139_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_139_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_139_BYTE_OFFSET = 13'h0958;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_139_ERR_INTRO_Q0_1_139_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_139_ERR_INTRO_Q0_1_139_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_139_ERR_INTRO_Q0_1_139_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_140_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_140_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_140_BYTE_OFFSET = 13'h095c;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_140_ERR_INTRO_Q0_1_140_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_140_ERR_INTRO_Q0_1_140_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_140_ERR_INTRO_Q0_1_140_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_141_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_141_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_141_BYTE_OFFSET = 13'h0960;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_141_ERR_INTRO_Q0_1_141_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_141_ERR_INTRO_Q0_1_141_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_141_ERR_INTRO_Q0_1_141_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_142_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_142_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_142_BYTE_OFFSET = 13'h0964;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_142_ERR_INTRO_Q0_1_142_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_142_ERR_INTRO_Q0_1_142_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_142_ERR_INTRO_Q0_1_142_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_143_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_143_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_143_BYTE_OFFSET = 13'h0968;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_143_ERR_INTRO_Q0_1_143_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_143_ERR_INTRO_Q0_1_143_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_143_ERR_INTRO_Q0_1_143_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_144_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_144_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_144_BYTE_OFFSET = 13'h096c;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_144_ERR_INTRO_Q0_1_144_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_144_ERR_INTRO_Q0_1_144_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_144_ERR_INTRO_Q0_1_144_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_145_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_145_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_145_BYTE_OFFSET = 13'h0970;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_145_ERR_INTRO_Q0_1_145_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_145_ERR_INTRO_Q0_1_145_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_145_ERR_INTRO_Q0_1_145_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_146_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_146_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_146_BYTE_OFFSET = 13'h0974;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_146_ERR_INTRO_Q0_1_146_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_146_ERR_INTRO_Q0_1_146_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_146_ERR_INTRO_Q0_1_146_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_147_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_147_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_147_BYTE_OFFSET = 13'h0978;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_147_ERR_INTRO_Q0_1_147_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_147_ERR_INTRO_Q0_1_147_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_147_ERR_INTRO_Q0_1_147_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_148_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_148_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_148_BYTE_OFFSET = 13'h097c;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_148_ERR_INTRO_Q0_1_148_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_148_ERR_INTRO_Q0_1_148_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_148_ERR_INTRO_Q0_1_148_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_149_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_149_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_149_BYTE_OFFSET = 13'h0980;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_149_ERR_INTRO_Q0_1_149_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_149_ERR_INTRO_Q0_1_149_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_149_ERR_INTRO_Q0_1_149_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_150_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_150_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_150_BYTE_OFFSET = 13'h0984;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_150_ERR_INTRO_Q0_1_150_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_150_ERR_INTRO_Q0_1_150_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_150_ERR_INTRO_Q0_1_150_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_151_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_151_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_151_BYTE_OFFSET = 13'h0988;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_151_ERR_INTRO_Q0_1_151_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_151_ERR_INTRO_Q0_1_151_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_151_ERR_INTRO_Q0_1_151_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_152_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_152_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_152_BYTE_OFFSET = 13'h098c;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_152_ERR_INTRO_Q0_1_152_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_152_ERR_INTRO_Q0_1_152_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_152_ERR_INTRO_Q0_1_152_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_153_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_153_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_153_BYTE_OFFSET = 13'h0990;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_153_ERR_INTRO_Q0_1_153_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_153_ERR_INTRO_Q0_1_153_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_153_ERR_INTRO_Q0_1_153_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_154_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_154_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_154_BYTE_OFFSET = 13'h0994;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_154_ERR_INTRO_Q0_1_154_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_154_ERR_INTRO_Q0_1_154_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_154_ERR_INTRO_Q0_1_154_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_155_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_155_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_155_BYTE_OFFSET = 13'h0998;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_155_ERR_INTRO_Q0_1_155_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_155_ERR_INTRO_Q0_1_155_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_155_ERR_INTRO_Q0_1_155_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_156_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_156_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_156_BYTE_OFFSET = 13'h099c;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_156_ERR_INTRO_Q0_1_156_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_156_ERR_INTRO_Q0_1_156_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_156_ERR_INTRO_Q0_1_156_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_157_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_157_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_157_BYTE_OFFSET = 13'h09a0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_157_ERR_INTRO_Q0_1_157_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_157_ERR_INTRO_Q0_1_157_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_157_ERR_INTRO_Q0_1_157_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_158_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_158_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_158_BYTE_OFFSET = 13'h09a4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_158_ERR_INTRO_Q0_1_158_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_158_ERR_INTRO_Q0_1_158_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_158_ERR_INTRO_Q0_1_158_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_159_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_159_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_159_BYTE_OFFSET = 13'h09a8;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_159_ERR_INTRO_Q0_1_159_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_159_ERR_INTRO_Q0_1_159_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_159_ERR_INTRO_Q0_1_159_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_160_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_160_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_160_BYTE_OFFSET = 13'h09ac;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_160_ERR_INTRO_Q0_1_160_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_160_ERR_INTRO_Q0_1_160_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_160_ERR_INTRO_Q0_1_160_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_161_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_161_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_161_BYTE_OFFSET = 13'h09b0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_161_ERR_INTRO_Q0_1_161_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_161_ERR_INTRO_Q0_1_161_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_161_ERR_INTRO_Q0_1_161_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_162_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_162_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_162_BYTE_OFFSET = 13'h09b4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_162_ERR_INTRO_Q0_1_162_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_162_ERR_INTRO_Q0_1_162_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_162_ERR_INTRO_Q0_1_162_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_163_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_163_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_163_BYTE_OFFSET = 13'h09b8;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_163_ERR_INTRO_Q0_1_163_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_163_ERR_INTRO_Q0_1_163_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_163_ERR_INTRO_Q0_1_163_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_164_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_164_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_164_BYTE_OFFSET = 13'h09bc;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_164_ERR_INTRO_Q0_1_164_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_164_ERR_INTRO_Q0_1_164_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_164_ERR_INTRO_Q0_1_164_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_165_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_165_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_165_BYTE_OFFSET = 13'h09c0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_165_ERR_INTRO_Q0_1_165_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_165_ERR_INTRO_Q0_1_165_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_165_ERR_INTRO_Q0_1_165_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_166_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_166_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_166_BYTE_OFFSET = 13'h09c4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_166_ERR_INTRO_Q0_1_166_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_166_ERR_INTRO_Q0_1_166_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_166_ERR_INTRO_Q0_1_166_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_167_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_167_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_167_BYTE_OFFSET = 13'h09c8;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_167_ERR_INTRO_Q0_1_167_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_167_ERR_INTRO_Q0_1_167_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_167_ERR_INTRO_Q0_1_167_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_168_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_168_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_168_BYTE_OFFSET = 13'h09cc;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_168_ERR_INTRO_Q0_1_168_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_168_ERR_INTRO_Q0_1_168_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_168_ERR_INTRO_Q0_1_168_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_169_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_169_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_169_BYTE_OFFSET = 13'h09d0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_169_ERR_INTRO_Q0_1_169_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_169_ERR_INTRO_Q0_1_169_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_169_ERR_INTRO_Q0_1_169_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_170_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_170_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_170_BYTE_OFFSET = 13'h09d4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_170_ERR_INTRO_Q0_1_170_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_170_ERR_INTRO_Q0_1_170_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_170_ERR_INTRO_Q0_1_170_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_171_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_171_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_171_BYTE_OFFSET = 13'h09d8;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_171_ERR_INTRO_Q0_1_171_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_171_ERR_INTRO_Q0_1_171_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_171_ERR_INTRO_Q0_1_171_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_172_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_172_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_172_BYTE_OFFSET = 13'h09dc;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_172_ERR_INTRO_Q0_1_172_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_172_ERR_INTRO_Q0_1_172_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_172_ERR_INTRO_Q0_1_172_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_173_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_173_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_173_BYTE_OFFSET = 13'h09e0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_173_ERR_INTRO_Q0_1_173_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_173_ERR_INTRO_Q0_1_173_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_173_ERR_INTRO_Q0_1_173_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_174_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_174_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_174_BYTE_OFFSET = 13'h09e4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_174_ERR_INTRO_Q0_1_174_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_174_ERR_INTRO_Q0_1_174_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_174_ERR_INTRO_Q0_1_174_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_175_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_175_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_175_BYTE_OFFSET = 13'h09e8;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_175_ERR_INTRO_Q0_1_175_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_175_ERR_INTRO_Q0_1_175_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_175_ERR_INTRO_Q0_1_175_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_176_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_176_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_176_BYTE_OFFSET = 13'h09ec;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_176_ERR_INTRO_Q0_1_176_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_176_ERR_INTRO_Q0_1_176_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_176_ERR_INTRO_Q0_1_176_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_177_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_177_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_177_BYTE_OFFSET = 13'h09f0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_177_ERR_INTRO_Q0_1_177_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_177_ERR_INTRO_Q0_1_177_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_177_ERR_INTRO_Q0_1_177_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_178_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_178_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_178_BYTE_OFFSET = 13'h09f4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_178_ERR_INTRO_Q0_1_178_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_178_ERR_INTRO_Q0_1_178_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_178_ERR_INTRO_Q0_1_178_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_179_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_179_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_179_BYTE_OFFSET = 13'h09f8;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_179_ERR_INTRO_Q0_1_179_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_179_ERR_INTRO_Q0_1_179_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_179_ERR_INTRO_Q0_1_179_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_180_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_180_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_180_BYTE_OFFSET = 13'h09fc;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_180_ERR_INTRO_Q0_1_180_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_180_ERR_INTRO_Q0_1_180_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_180_ERR_INTRO_Q0_1_180_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_181_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_181_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_181_BYTE_OFFSET = 13'h0a00;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_181_ERR_INTRO_Q0_1_181_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_181_ERR_INTRO_Q0_1_181_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_181_ERR_INTRO_Q0_1_181_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_182_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_182_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_182_BYTE_OFFSET = 13'h0a04;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_182_ERR_INTRO_Q0_1_182_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_182_ERR_INTRO_Q0_1_182_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_182_ERR_INTRO_Q0_1_182_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_183_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_183_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_183_BYTE_OFFSET = 13'h0a08;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_183_ERR_INTRO_Q0_1_183_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_183_ERR_INTRO_Q0_1_183_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_183_ERR_INTRO_Q0_1_183_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_184_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_184_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_184_BYTE_OFFSET = 13'h0a0c;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_184_ERR_INTRO_Q0_1_184_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_184_ERR_INTRO_Q0_1_184_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_184_ERR_INTRO_Q0_1_184_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_185_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_185_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_185_BYTE_OFFSET = 13'h0a10;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_185_ERR_INTRO_Q0_1_185_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_185_ERR_INTRO_Q0_1_185_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_185_ERR_INTRO_Q0_1_185_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_186_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_186_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_186_BYTE_OFFSET = 13'h0a14;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_186_ERR_INTRO_Q0_1_186_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_186_ERR_INTRO_Q0_1_186_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_186_ERR_INTRO_Q0_1_186_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_187_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_187_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_187_BYTE_OFFSET = 13'h0a18;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_187_ERR_INTRO_Q0_1_187_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_187_ERR_INTRO_Q0_1_187_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_187_ERR_INTRO_Q0_1_187_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_188_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_188_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_188_BYTE_OFFSET = 13'h0a1c;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_188_ERR_INTRO_Q0_1_188_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_188_ERR_INTRO_Q0_1_188_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_188_ERR_INTRO_Q0_1_188_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_189_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_189_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_189_BYTE_OFFSET = 13'h0a20;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_189_ERR_INTRO_Q0_1_189_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_189_ERR_INTRO_Q0_1_189_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_189_ERR_INTRO_Q0_1_189_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_190_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_190_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_190_BYTE_OFFSET = 13'h0a24;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_190_ERR_INTRO_Q0_1_190_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_190_ERR_INTRO_Q0_1_190_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_190_ERR_INTRO_Q0_1_190_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_191_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_191_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_191_BYTE_OFFSET = 13'h0a28;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_191_ERR_INTRO_Q0_1_191_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_191_ERR_INTRO_Q0_1_191_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_191_ERR_INTRO_Q0_1_191_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_192_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_192_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_192_BYTE_OFFSET = 13'h0a2c;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_192_ERR_INTRO_Q0_1_192_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_192_ERR_INTRO_Q0_1_192_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_192_ERR_INTRO_Q0_1_192_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_193_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_193_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_193_BYTE_OFFSET = 13'h0a30;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_193_ERR_INTRO_Q0_1_193_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_193_ERR_INTRO_Q0_1_193_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_193_ERR_INTRO_Q0_1_193_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_194_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_194_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_194_BYTE_OFFSET = 13'h0a34;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_194_ERR_INTRO_Q0_1_194_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_194_ERR_INTRO_Q0_1_194_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_194_ERR_INTRO_Q0_1_194_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_195_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_195_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_195_BYTE_OFFSET = 13'h0a38;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_195_ERR_INTRO_Q0_1_195_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_195_ERR_INTRO_Q0_1_195_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_195_ERR_INTRO_Q0_1_195_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_196_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_196_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_196_BYTE_OFFSET = 13'h0a3c;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_196_ERR_INTRO_Q0_1_196_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_196_ERR_INTRO_Q0_1_196_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_196_ERR_INTRO_Q0_1_196_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_197_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_197_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_197_BYTE_OFFSET = 13'h0a40;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_197_ERR_INTRO_Q0_1_197_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_197_ERR_INTRO_Q0_1_197_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_197_ERR_INTRO_Q0_1_197_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_198_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_198_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_198_BYTE_OFFSET = 13'h0a44;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_198_ERR_INTRO_Q0_1_198_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_198_ERR_INTRO_Q0_1_198_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_198_ERR_INTRO_Q0_1_198_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_199_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_199_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_199_BYTE_OFFSET = 13'h0a48;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_199_ERR_INTRO_Q0_1_199_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_199_ERR_INTRO_Q0_1_199_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_199_ERR_INTRO_Q0_1_199_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_200_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_200_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_200_BYTE_OFFSET = 13'h0a4c;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_200_ERR_INTRO_Q0_1_200_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_200_ERR_INTRO_Q0_1_200_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_200_ERR_INTRO_Q0_1_200_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_201_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_201_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_201_BYTE_OFFSET = 13'h0a50;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_201_ERR_INTRO_Q0_1_201_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_201_ERR_INTRO_Q0_1_201_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_201_ERR_INTRO_Q0_1_201_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_202_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_202_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_202_BYTE_OFFSET = 13'h0a54;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_202_ERR_INTRO_Q0_1_202_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_202_ERR_INTRO_Q0_1_202_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_202_ERR_INTRO_Q0_1_202_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_203_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_203_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_203_BYTE_OFFSET = 13'h0a58;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_203_ERR_INTRO_Q0_1_203_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_203_ERR_INTRO_Q0_1_203_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_203_ERR_INTRO_Q0_1_203_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_204_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_204_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_204_BYTE_OFFSET = 13'h0a5c;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_204_ERR_INTRO_Q0_1_204_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_204_ERR_INTRO_Q0_1_204_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_204_ERR_INTRO_Q0_1_204_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_205_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_205_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_205_BYTE_OFFSET = 13'h0a60;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_205_ERR_INTRO_Q0_1_205_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_205_ERR_INTRO_Q0_1_205_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_205_ERR_INTRO_Q0_1_205_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_206_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_206_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_206_BYTE_OFFSET = 13'h0a64;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_206_ERR_INTRO_Q0_1_206_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_206_ERR_INTRO_Q0_1_206_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_206_ERR_INTRO_Q0_1_206_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_207_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_207_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_Q0_1_INTRO_207_BYTE_OFFSET = 13'h0a68;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_207_ERR_INTRO_Q0_1_207_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_Q0_1_INTRO_207_ERR_INTRO_Q0_1_207_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_Q0_1_INTRO_207_ERR_INTRO_Q0_1_207_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_0_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_0_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_0_BYTE_OFFSET = 13'h0a6c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_0_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_0_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_0_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_1_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_1_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_1_BYTE_OFFSET = 13'h0a70;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_1_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_1_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_1_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_2_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_2_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_2_BYTE_OFFSET = 13'h0a74;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_2_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_2_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_2_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_3_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_3_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_3_BYTE_OFFSET = 13'h0a78;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_3_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_3_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_3_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_4_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_4_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_4_BYTE_OFFSET = 13'h0a7c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_4_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_4_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_4_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_5_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_5_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_5_BYTE_OFFSET = 13'h0a80;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_5_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_5_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_5_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_6_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_6_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_6_BYTE_OFFSET = 13'h0a84;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_6_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_6_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_6_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_7_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_7_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_7_BYTE_OFFSET = 13'h0a88;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_7_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_7_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_7_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_8_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_8_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_8_BYTE_OFFSET = 13'h0a8c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_8_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_8_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_8_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_9_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_9_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_9_BYTE_OFFSET = 13'h0a90;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_9_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_9_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_9_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_10_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_10_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_10_BYTE_OFFSET = 13'h0a94;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_10_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_10_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_10_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_11_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_11_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_11_BYTE_OFFSET = 13'h0a98;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_11_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_11_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_11_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_12_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_12_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_12_BYTE_OFFSET = 13'h0a9c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_12_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_12_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_12_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_13_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_13_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_13_BYTE_OFFSET = 13'h0aa0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_13_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_13_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_13_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_14_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_14_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_14_BYTE_OFFSET = 13'h0aa4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_14_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_14_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_14_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_15_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_15_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_15_BYTE_OFFSET = 13'h0aa8;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_15_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_15_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_15_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_16_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_16_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_16_BYTE_OFFSET = 13'h0aac;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_16_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_16_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_16_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_17_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_17_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_17_BYTE_OFFSET = 13'h0ab0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_17_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_17_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_17_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_18_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_18_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_18_BYTE_OFFSET = 13'h0ab4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_18_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_18_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_18_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_19_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_19_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_19_BYTE_OFFSET = 13'h0ab8;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_19_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_19_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_19_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_20_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_20_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_20_BYTE_OFFSET = 13'h0abc;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_20_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_20_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_20_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_21_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_21_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_21_BYTE_OFFSET = 13'h0ac0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_21_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_21_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_21_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_22_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_22_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_22_BYTE_OFFSET = 13'h0ac4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_22_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_22_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_22_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_23_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_23_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_23_BYTE_OFFSET = 13'h0ac8;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_23_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_23_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_23_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_24_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_24_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_24_BYTE_OFFSET = 13'h0acc;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_24_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_24_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_24_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_25_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_25_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_25_BYTE_OFFSET = 13'h0ad0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_25_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_25_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_25_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_26_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_26_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_26_BYTE_OFFSET = 13'h0ad4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_26_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_26_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_26_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_27_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_27_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_27_BYTE_OFFSET = 13'h0ad8;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_27_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_27_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_27_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_28_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_28_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_28_BYTE_OFFSET = 13'h0adc;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_28_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_28_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_28_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_29_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_29_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_29_BYTE_OFFSET = 13'h0ae0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_29_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_29_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_29_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_30_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_30_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_30_BYTE_OFFSET = 13'h0ae4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_30_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_30_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_30_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_31_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_31_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_31_BYTE_OFFSET = 13'h0ae8;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_31_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_31_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_31_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_32_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_32_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_32_BYTE_OFFSET = 13'h0aec;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_32_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_32_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_32_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_33_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_33_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_33_BYTE_OFFSET = 13'h0af0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_33_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_33_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_33_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_34_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_34_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_34_BYTE_OFFSET = 13'h0af4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_34_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_34_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_34_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_35_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_35_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_35_BYTE_OFFSET = 13'h0af8;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_35_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_35_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_35_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_36_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_36_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_36_BYTE_OFFSET = 13'h0afc;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_36_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_36_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_36_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_37_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_37_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_37_BYTE_OFFSET = 13'h0b00;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_37_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_37_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_37_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_38_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_38_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_38_BYTE_OFFSET = 13'h0b04;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_38_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_38_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_38_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_39_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_39_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_39_BYTE_OFFSET = 13'h0b08;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_39_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_39_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_39_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_40_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_40_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_40_BYTE_OFFSET = 13'h0b0c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_40_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_40_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_40_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_41_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_41_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_41_BYTE_OFFSET = 13'h0b10;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_41_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_41_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_41_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_42_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_42_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_42_BYTE_OFFSET = 13'h0b14;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_42_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_42_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_42_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_43_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_43_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_43_BYTE_OFFSET = 13'h0b18;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_43_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_43_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_43_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_44_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_44_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_44_BYTE_OFFSET = 13'h0b1c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_44_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_44_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_44_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_45_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_45_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_45_BYTE_OFFSET = 13'h0b20;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_45_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_45_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_45_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_46_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_46_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_46_BYTE_OFFSET = 13'h0b24;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_46_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_46_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_46_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_47_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_47_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_47_BYTE_OFFSET = 13'h0b28;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_47_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_47_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_47_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_48_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_48_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_48_BYTE_OFFSET = 13'h0b2c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_48_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_48_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_48_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_49_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_49_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_49_BYTE_OFFSET = 13'h0b30;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_49_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_49_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_49_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_50_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_50_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_50_BYTE_OFFSET = 13'h0b34;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_50_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_50_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_50_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_51_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_51_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_51_BYTE_OFFSET = 13'h0b38;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_51_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_51_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_51_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_52_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_52_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_52_BYTE_OFFSET = 13'h0b3c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_52_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_52_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_52_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_53_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_53_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_53_BYTE_OFFSET = 13'h0b40;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_53_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_53_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_53_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_54_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_54_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_54_BYTE_OFFSET = 13'h0b44;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_54_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_54_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_54_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_55_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_55_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_55_BYTE_OFFSET = 13'h0b48;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_55_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_55_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_55_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_56_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_56_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_56_BYTE_OFFSET = 13'h0b4c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_56_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_56_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_56_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_57_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_57_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_57_BYTE_OFFSET = 13'h0b50;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_57_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_57_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_57_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_58_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_58_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_58_BYTE_OFFSET = 13'h0b54;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_58_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_58_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_58_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_59_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_59_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_59_BYTE_OFFSET = 13'h0b58;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_59_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_59_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_59_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_60_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_60_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_60_BYTE_OFFSET = 13'h0b5c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_60_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_60_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_60_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_61_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_61_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_61_BYTE_OFFSET = 13'h0b60;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_61_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_61_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_61_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_62_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_62_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_62_BYTE_OFFSET = 13'h0b64;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_62_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_62_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_62_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_63_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_63_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_63_BYTE_OFFSET = 13'h0b68;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_63_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_63_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_63_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_64_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_64_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_64_BYTE_OFFSET = 13'h0b6c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_64_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_64_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_64_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_65_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_65_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_65_BYTE_OFFSET = 13'h0b70;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_65_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_65_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_65_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_66_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_66_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_66_BYTE_OFFSET = 13'h0b74;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_66_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_66_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_66_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_67_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_67_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_67_BYTE_OFFSET = 13'h0b78;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_67_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_67_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_67_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_68_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_68_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_68_BYTE_OFFSET = 13'h0b7c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_68_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_68_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_68_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_69_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_69_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_69_BYTE_OFFSET = 13'h0b80;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_69_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_69_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_69_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_70_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_70_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_70_BYTE_OFFSET = 13'h0b84;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_70_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_70_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_70_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_71_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_71_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_71_BYTE_OFFSET = 13'h0b88;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_71_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_71_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_71_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_72_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_72_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_72_BYTE_OFFSET = 13'h0b8c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_72_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_72_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_72_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_73_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_73_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_73_BYTE_OFFSET = 13'h0b90;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_73_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_73_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_73_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_74_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_74_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_74_BYTE_OFFSET = 13'h0b94;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_74_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_74_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_74_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_75_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_75_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_75_BYTE_OFFSET = 13'h0b98;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_75_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_75_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_75_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_76_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_76_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_76_BYTE_OFFSET = 13'h0b9c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_76_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_76_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_76_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_77_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_77_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_77_BYTE_OFFSET = 13'h0ba0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_77_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_77_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_77_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_78_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_78_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_78_BYTE_OFFSET = 13'h0ba4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_78_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_78_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_78_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_79_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_79_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_79_BYTE_OFFSET = 13'h0ba8;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_79_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_79_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_79_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_80_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_80_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_80_BYTE_OFFSET = 13'h0bac;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_80_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_80_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_80_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_81_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_81_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_81_BYTE_OFFSET = 13'h0bb0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_81_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_81_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_81_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_82_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_82_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_82_BYTE_OFFSET = 13'h0bb4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_82_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_82_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_82_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_83_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_83_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_83_BYTE_OFFSET = 13'h0bb8;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_83_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_83_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_83_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_84_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_84_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_84_BYTE_OFFSET = 13'h0bbc;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_84_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_84_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_84_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_85_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_85_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_85_BYTE_OFFSET = 13'h0bc0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_85_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_85_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_85_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_86_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_86_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_86_BYTE_OFFSET = 13'h0bc4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_86_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_86_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_86_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_87_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_87_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_87_BYTE_OFFSET = 13'h0bc8;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_87_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_87_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_87_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_88_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_88_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_88_BYTE_OFFSET = 13'h0bcc;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_88_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_88_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_88_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_89_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_89_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_89_BYTE_OFFSET = 13'h0bd0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_89_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_89_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_89_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_90_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_90_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_90_BYTE_OFFSET = 13'h0bd4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_90_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_90_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_90_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_91_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_91_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_91_BYTE_OFFSET = 13'h0bd8;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_91_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_91_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_91_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_92_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_92_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_92_BYTE_OFFSET = 13'h0bdc;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_92_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_92_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_92_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_93_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_93_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_93_BYTE_OFFSET = 13'h0be0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_93_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_93_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_93_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_94_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_94_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_94_BYTE_OFFSET = 13'h0be4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_94_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_94_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_94_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_95_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_95_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_95_BYTE_OFFSET = 13'h0be8;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_95_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_95_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_95_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_96_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_96_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_96_BYTE_OFFSET = 13'h0bec;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_96_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_96_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_96_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_97_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_97_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_97_BYTE_OFFSET = 13'h0bf0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_97_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_97_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_97_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_98_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_98_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_98_BYTE_OFFSET = 13'h0bf4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_98_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_98_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_98_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_99_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_99_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_99_BYTE_OFFSET = 13'h0bf8;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_99_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_99_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_99_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_100_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_100_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_100_BYTE_OFFSET = 13'h0bfc;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_100_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_100_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_100_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_101_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_101_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_101_BYTE_OFFSET = 13'h0c00;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_101_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_101_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_101_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_102_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_102_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_102_BYTE_OFFSET = 13'h0c04;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_102_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_102_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_102_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_103_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_103_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_103_BYTE_OFFSET = 13'h0c08;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_103_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_103_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_103_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_104_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_104_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_104_BYTE_OFFSET = 13'h0c0c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_104_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_104_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_104_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_105_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_105_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_105_BYTE_OFFSET = 13'h0c10;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_105_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_105_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_105_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_106_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_106_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_106_BYTE_OFFSET = 13'h0c14;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_106_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_106_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_106_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_107_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_107_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_107_BYTE_OFFSET = 13'h0c18;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_107_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_107_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_107_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_108_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_108_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_108_BYTE_OFFSET = 13'h0c1c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_108_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_108_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_108_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_109_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_109_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_109_BYTE_OFFSET = 13'h0c20;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_109_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_109_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_109_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_110_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_110_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_110_BYTE_OFFSET = 13'h0c24;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_110_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_110_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_110_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_111_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_111_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_111_BYTE_OFFSET = 13'h0c28;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_111_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_111_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_111_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_112_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_112_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_112_BYTE_OFFSET = 13'h0c2c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_112_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_112_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_112_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_113_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_113_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_113_BYTE_OFFSET = 13'h0c30;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_113_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_113_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_113_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_114_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_114_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_114_BYTE_OFFSET = 13'h0c34;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_114_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_114_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_114_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_115_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_115_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_115_BYTE_OFFSET = 13'h0c38;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_115_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_115_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_115_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_116_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_116_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_116_BYTE_OFFSET = 13'h0c3c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_116_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_116_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_116_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_117_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_117_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_117_BYTE_OFFSET = 13'h0c40;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_117_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_117_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_117_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_118_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_118_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_118_BYTE_OFFSET = 13'h0c44;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_118_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_118_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_118_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_119_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_119_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_119_BYTE_OFFSET = 13'h0c48;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_119_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_119_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_119_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_120_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_120_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_120_BYTE_OFFSET = 13'h0c4c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_120_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_120_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_120_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_121_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_121_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_121_BYTE_OFFSET = 13'h0c50;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_121_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_121_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_121_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_122_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_122_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_122_BYTE_OFFSET = 13'h0c54;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_122_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_122_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_122_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_123_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_123_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_123_BYTE_OFFSET = 13'h0c58;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_123_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_123_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_123_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_124_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_124_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_124_BYTE_OFFSET = 13'h0c5c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_124_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_124_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_124_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_125_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_125_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_125_BYTE_OFFSET = 13'h0c60;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_125_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_125_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_125_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_126_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_126_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_126_BYTE_OFFSET = 13'h0c64;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_126_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_126_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_126_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_127_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_127_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_127_BYTE_OFFSET = 13'h0c68;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_127_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_127_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_127_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_128_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_128_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_128_BYTE_OFFSET = 13'h0c6c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_128_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_128_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_128_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_129_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_129_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_129_BYTE_OFFSET = 13'h0c70;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_129_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_129_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_129_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_130_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_130_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_130_BYTE_OFFSET = 13'h0c74;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_130_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_130_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_130_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_131_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_131_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_131_BYTE_OFFSET = 13'h0c78;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_131_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_131_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_131_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_132_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_132_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_132_BYTE_OFFSET = 13'h0c7c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_132_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_132_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_132_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_133_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_133_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_133_BYTE_OFFSET = 13'h0c80;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_133_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_133_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_133_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_134_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_134_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_134_BYTE_OFFSET = 13'h0c84;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_134_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_134_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_134_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_135_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_135_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_135_BYTE_OFFSET = 13'h0c88;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_135_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_135_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_135_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_136_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_136_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_136_BYTE_OFFSET = 13'h0c8c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_136_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_136_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_136_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_137_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_137_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_137_BYTE_OFFSET = 13'h0c90;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_137_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_137_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_137_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_138_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_138_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_138_BYTE_OFFSET = 13'h0c94;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_138_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_138_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_138_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_139_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_139_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_139_BYTE_OFFSET = 13'h0c98;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_139_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_139_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_139_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_140_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_140_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_140_BYTE_OFFSET = 13'h0c9c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_140_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_140_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_140_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_141_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_141_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_141_BYTE_OFFSET = 13'h0ca0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_141_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_141_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_141_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_142_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_142_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_142_BYTE_OFFSET = 13'h0ca4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_142_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_142_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_142_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_143_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_143_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_143_BYTE_OFFSET = 13'h0ca8;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_143_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_143_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_143_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_144_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_144_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_144_BYTE_OFFSET = 13'h0cac;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_144_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_144_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_144_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_145_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_145_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_145_BYTE_OFFSET = 13'h0cb0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_145_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_145_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_145_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_146_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_146_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_146_BYTE_OFFSET = 13'h0cb4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_146_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_146_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_146_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_147_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_147_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_147_BYTE_OFFSET = 13'h0cb8;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_147_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_147_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_147_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_148_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_148_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_148_BYTE_OFFSET = 13'h0cbc;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_148_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_148_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_148_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_149_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_149_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_149_BYTE_OFFSET = 13'h0cc0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_149_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_149_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_149_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_150_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_150_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_150_BYTE_OFFSET = 13'h0cc4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_150_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_150_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_150_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_151_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_151_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_151_BYTE_OFFSET = 13'h0cc8;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_151_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_151_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_151_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_152_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_152_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_152_BYTE_OFFSET = 13'h0ccc;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_152_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_152_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_152_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_153_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_153_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_153_BYTE_OFFSET = 13'h0cd0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_153_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_153_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_153_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_154_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_154_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_154_BYTE_OFFSET = 13'h0cd4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_154_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_154_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_154_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_155_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_155_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_155_BYTE_OFFSET = 13'h0cd8;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_155_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_155_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_155_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_156_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_156_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_156_BYTE_OFFSET = 13'h0cdc;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_156_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_156_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_156_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_157_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_157_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_157_BYTE_OFFSET = 13'h0ce0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_157_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_157_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_157_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_158_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_158_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_158_BYTE_OFFSET = 13'h0ce4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_158_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_158_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_158_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_159_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_159_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_159_BYTE_OFFSET = 13'h0ce8;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_159_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_159_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_159_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_160_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_160_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_160_BYTE_OFFSET = 13'h0cec;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_160_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_160_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_160_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_161_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_161_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_161_BYTE_OFFSET = 13'h0cf0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_161_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_161_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_161_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_162_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_162_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_162_BYTE_OFFSET = 13'h0cf4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_162_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_162_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_162_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_163_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_163_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_163_BYTE_OFFSET = 13'h0cf8;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_163_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_163_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_163_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_164_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_164_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_164_BYTE_OFFSET = 13'h0cfc;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_164_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_164_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_164_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_165_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_165_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_165_BYTE_OFFSET = 13'h0d00;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_165_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_165_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_165_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_166_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_166_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_166_BYTE_OFFSET = 13'h0d04;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_166_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_166_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_166_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_167_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_167_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_167_BYTE_OFFSET = 13'h0d08;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_167_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_167_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_167_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_168_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_168_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_168_BYTE_OFFSET = 13'h0d0c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_168_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_168_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_168_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_169_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_169_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_169_BYTE_OFFSET = 13'h0d10;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_169_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_169_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_169_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_170_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_170_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_170_BYTE_OFFSET = 13'h0d14;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_170_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_170_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_170_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_171_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_171_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_171_BYTE_OFFSET = 13'h0d18;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_171_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_171_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_171_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_172_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_172_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_172_BYTE_OFFSET = 13'h0d1c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_172_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_172_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_172_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_173_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_173_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_173_BYTE_OFFSET = 13'h0d20;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_173_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_173_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_173_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_174_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_174_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_174_BYTE_OFFSET = 13'h0d24;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_174_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_174_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_174_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_175_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_175_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_175_BYTE_OFFSET = 13'h0d28;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_175_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_175_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_175_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_176_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_176_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_176_BYTE_OFFSET = 13'h0d2c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_176_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_176_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_176_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_177_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_177_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_177_BYTE_OFFSET = 13'h0d30;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_177_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_177_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_177_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_178_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_178_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_178_BYTE_OFFSET = 13'h0d34;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_178_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_178_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_178_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_179_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_179_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_179_BYTE_OFFSET = 13'h0d38;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_179_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_179_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_179_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_180_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_180_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_180_BYTE_OFFSET = 13'h0d3c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_180_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_180_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_180_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_181_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_181_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_181_BYTE_OFFSET = 13'h0d40;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_181_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_181_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_181_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_182_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_182_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_182_BYTE_OFFSET = 13'h0d44;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_182_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_182_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_182_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_183_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_183_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_183_BYTE_OFFSET = 13'h0d48;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_183_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_183_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_183_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_184_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_184_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_184_BYTE_OFFSET = 13'h0d4c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_184_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_184_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_184_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_185_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_185_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_185_BYTE_OFFSET = 13'h0d50;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_185_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_185_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_185_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_186_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_186_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_186_BYTE_OFFSET = 13'h0d54;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_186_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_186_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_186_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_187_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_187_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_187_BYTE_OFFSET = 13'h0d58;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_187_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_187_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_187_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_188_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_188_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_188_BYTE_OFFSET = 13'h0d5c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_188_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_188_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_188_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_189_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_189_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_189_BYTE_OFFSET = 13'h0d60;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_189_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_189_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_189_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_190_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_190_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_190_BYTE_OFFSET = 13'h0d64;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_190_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_190_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_190_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_191_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_191_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_191_BYTE_OFFSET = 13'h0d68;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_191_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_191_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_191_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_192_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_192_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_192_BYTE_OFFSET = 13'h0d6c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_192_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_192_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_192_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_193_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_193_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_193_BYTE_OFFSET = 13'h0d70;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_193_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_193_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_193_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_194_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_194_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_194_BYTE_OFFSET = 13'h0d74;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_194_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_194_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_194_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_195_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_195_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_195_BYTE_OFFSET = 13'h0d78;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_195_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_195_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_195_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_196_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_196_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_196_BYTE_OFFSET = 13'h0d7c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_196_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_196_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_196_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_197_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_197_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_197_BYTE_OFFSET = 13'h0d80;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_197_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_197_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_197_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_198_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_198_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_198_BYTE_OFFSET = 13'h0d84;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_198_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_198_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_198_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_199_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_199_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_199_BYTE_OFFSET = 13'h0d88;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_199_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_199_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_199_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_200_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_200_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_200_BYTE_OFFSET = 13'h0d8c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_200_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_200_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_200_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_201_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_201_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_201_BYTE_OFFSET = 13'h0d90;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_201_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_201_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_201_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_202_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_202_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_202_BYTE_OFFSET = 13'h0d94;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_202_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_202_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_202_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_203_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_203_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_203_BYTE_OFFSET = 13'h0d98;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_203_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_203_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_203_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_204_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_204_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_204_BYTE_OFFSET = 13'h0d9c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_204_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_204_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_204_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_205_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_205_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_205_BYTE_OFFSET = 13'h0da0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_205_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_205_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_205_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_206_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_206_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_206_BYTE_OFFSET = 13'h0da4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_206_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_206_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_206_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_207_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_207_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_0_207_BYTE_OFFSET = 13'h0da8;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_207_CWORD_Q0_0_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_0_207_CWORD_Q0_0_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_0_207_CWORD_Q0_0_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_0_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_0_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_0_BYTE_OFFSET = 13'h0dac;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_0_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_0_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_0_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_1_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_1_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_1_BYTE_OFFSET = 13'h0db0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_1_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_1_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_1_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_2_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_2_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_2_BYTE_OFFSET = 13'h0db4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_2_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_2_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_2_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_3_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_3_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_3_BYTE_OFFSET = 13'h0db8;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_3_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_3_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_3_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_4_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_4_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_4_BYTE_OFFSET = 13'h0dbc;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_4_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_4_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_4_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_5_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_5_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_5_BYTE_OFFSET = 13'h0dc0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_5_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_5_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_5_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_6_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_6_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_6_BYTE_OFFSET = 13'h0dc4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_6_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_6_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_6_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_7_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_7_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_7_BYTE_OFFSET = 13'h0dc8;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_7_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_7_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_7_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_8_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_8_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_8_BYTE_OFFSET = 13'h0dcc;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_8_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_8_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_8_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_9_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_9_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_9_BYTE_OFFSET = 13'h0dd0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_9_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_9_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_9_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_10_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_10_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_10_BYTE_OFFSET = 13'h0dd4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_10_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_10_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_10_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_11_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_11_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_11_BYTE_OFFSET = 13'h0dd8;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_11_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_11_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_11_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_12_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_12_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_12_BYTE_OFFSET = 13'h0ddc;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_12_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_12_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_12_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_13_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_13_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_13_BYTE_OFFSET = 13'h0de0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_13_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_13_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_13_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_14_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_14_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_14_BYTE_OFFSET = 13'h0de4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_14_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_14_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_14_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_15_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_15_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_15_BYTE_OFFSET = 13'h0de8;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_15_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_15_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_15_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_16_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_16_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_16_BYTE_OFFSET = 13'h0dec;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_16_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_16_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_16_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_17_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_17_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_17_BYTE_OFFSET = 13'h0df0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_17_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_17_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_17_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_18_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_18_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_18_BYTE_OFFSET = 13'h0df4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_18_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_18_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_18_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_19_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_19_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_19_BYTE_OFFSET = 13'h0df8;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_19_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_19_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_19_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_20_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_20_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_20_BYTE_OFFSET = 13'h0dfc;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_20_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_20_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_20_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_21_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_21_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_21_BYTE_OFFSET = 13'h0e00;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_21_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_21_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_21_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_22_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_22_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_22_BYTE_OFFSET = 13'h0e04;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_22_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_22_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_22_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_23_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_23_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_23_BYTE_OFFSET = 13'h0e08;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_23_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_23_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_23_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_24_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_24_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_24_BYTE_OFFSET = 13'h0e0c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_24_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_24_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_24_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_25_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_25_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_25_BYTE_OFFSET = 13'h0e10;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_25_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_25_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_25_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_26_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_26_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_26_BYTE_OFFSET = 13'h0e14;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_26_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_26_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_26_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_27_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_27_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_27_BYTE_OFFSET = 13'h0e18;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_27_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_27_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_27_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_28_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_28_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_28_BYTE_OFFSET = 13'h0e1c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_28_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_28_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_28_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_29_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_29_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_29_BYTE_OFFSET = 13'h0e20;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_29_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_29_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_29_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_30_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_30_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_30_BYTE_OFFSET = 13'h0e24;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_30_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_30_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_30_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_31_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_31_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_31_BYTE_OFFSET = 13'h0e28;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_31_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_31_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_31_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_32_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_32_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_32_BYTE_OFFSET = 13'h0e2c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_32_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_32_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_32_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_33_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_33_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_33_BYTE_OFFSET = 13'h0e30;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_33_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_33_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_33_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_34_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_34_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_34_BYTE_OFFSET = 13'h0e34;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_34_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_34_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_34_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_35_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_35_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_35_BYTE_OFFSET = 13'h0e38;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_35_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_35_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_35_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_36_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_36_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_36_BYTE_OFFSET = 13'h0e3c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_36_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_36_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_36_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_37_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_37_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_37_BYTE_OFFSET = 13'h0e40;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_37_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_37_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_37_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_38_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_38_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_38_BYTE_OFFSET = 13'h0e44;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_38_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_38_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_38_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_39_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_39_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_39_BYTE_OFFSET = 13'h0e48;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_39_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_39_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_39_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_40_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_40_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_40_BYTE_OFFSET = 13'h0e4c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_40_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_40_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_40_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_41_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_41_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_41_BYTE_OFFSET = 13'h0e50;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_41_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_41_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_41_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_42_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_42_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_42_BYTE_OFFSET = 13'h0e54;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_42_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_42_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_42_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_43_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_43_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_43_BYTE_OFFSET = 13'h0e58;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_43_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_43_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_43_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_44_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_44_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_44_BYTE_OFFSET = 13'h0e5c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_44_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_44_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_44_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_45_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_45_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_45_BYTE_OFFSET = 13'h0e60;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_45_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_45_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_45_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_46_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_46_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_46_BYTE_OFFSET = 13'h0e64;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_46_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_46_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_46_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_47_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_47_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_47_BYTE_OFFSET = 13'h0e68;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_47_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_47_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_47_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_48_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_48_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_48_BYTE_OFFSET = 13'h0e6c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_48_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_48_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_48_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_49_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_49_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_49_BYTE_OFFSET = 13'h0e70;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_49_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_49_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_49_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_50_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_50_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_50_BYTE_OFFSET = 13'h0e74;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_50_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_50_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_50_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_51_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_51_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_51_BYTE_OFFSET = 13'h0e78;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_51_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_51_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_51_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_52_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_52_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_52_BYTE_OFFSET = 13'h0e7c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_52_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_52_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_52_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_53_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_53_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_53_BYTE_OFFSET = 13'h0e80;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_53_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_53_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_53_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_54_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_54_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_54_BYTE_OFFSET = 13'h0e84;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_54_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_54_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_54_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_55_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_55_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_55_BYTE_OFFSET = 13'h0e88;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_55_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_55_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_55_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_56_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_56_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_56_BYTE_OFFSET = 13'h0e8c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_56_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_56_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_56_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_57_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_57_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_57_BYTE_OFFSET = 13'h0e90;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_57_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_57_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_57_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_58_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_58_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_58_BYTE_OFFSET = 13'h0e94;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_58_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_58_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_58_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_59_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_59_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_59_BYTE_OFFSET = 13'h0e98;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_59_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_59_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_59_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_60_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_60_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_60_BYTE_OFFSET = 13'h0e9c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_60_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_60_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_60_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_61_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_61_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_61_BYTE_OFFSET = 13'h0ea0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_61_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_61_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_61_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_62_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_62_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_62_BYTE_OFFSET = 13'h0ea4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_62_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_62_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_62_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_63_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_63_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_63_BYTE_OFFSET = 13'h0ea8;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_63_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_63_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_63_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_64_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_64_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_64_BYTE_OFFSET = 13'h0eac;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_64_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_64_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_64_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_65_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_65_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_65_BYTE_OFFSET = 13'h0eb0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_65_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_65_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_65_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_66_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_66_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_66_BYTE_OFFSET = 13'h0eb4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_66_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_66_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_66_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_67_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_67_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_67_BYTE_OFFSET = 13'h0eb8;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_67_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_67_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_67_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_68_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_68_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_68_BYTE_OFFSET = 13'h0ebc;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_68_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_68_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_68_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_69_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_69_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_69_BYTE_OFFSET = 13'h0ec0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_69_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_69_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_69_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_70_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_70_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_70_BYTE_OFFSET = 13'h0ec4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_70_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_70_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_70_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_71_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_71_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_71_BYTE_OFFSET = 13'h0ec8;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_71_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_71_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_71_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_72_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_72_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_72_BYTE_OFFSET = 13'h0ecc;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_72_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_72_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_72_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_73_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_73_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_73_BYTE_OFFSET = 13'h0ed0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_73_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_73_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_73_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_74_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_74_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_74_BYTE_OFFSET = 13'h0ed4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_74_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_74_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_74_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_75_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_75_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_75_BYTE_OFFSET = 13'h0ed8;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_75_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_75_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_75_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_76_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_76_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_76_BYTE_OFFSET = 13'h0edc;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_76_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_76_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_76_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_77_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_77_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_77_BYTE_OFFSET = 13'h0ee0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_77_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_77_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_77_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_78_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_78_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_78_BYTE_OFFSET = 13'h0ee4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_78_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_78_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_78_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_79_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_79_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_79_BYTE_OFFSET = 13'h0ee8;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_79_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_79_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_79_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_80_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_80_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_80_BYTE_OFFSET = 13'h0eec;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_80_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_80_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_80_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_81_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_81_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_81_BYTE_OFFSET = 13'h0ef0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_81_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_81_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_81_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_82_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_82_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_82_BYTE_OFFSET = 13'h0ef4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_82_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_82_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_82_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_83_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_83_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_83_BYTE_OFFSET = 13'h0ef8;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_83_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_83_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_83_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_84_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_84_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_84_BYTE_OFFSET = 13'h0efc;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_84_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_84_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_84_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_85_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_85_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_85_BYTE_OFFSET = 13'h0f00;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_85_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_85_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_85_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_86_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_86_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_86_BYTE_OFFSET = 13'h0f04;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_86_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_86_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_86_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_87_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_87_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_87_BYTE_OFFSET = 13'h0f08;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_87_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_87_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_87_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_88_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_88_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_88_BYTE_OFFSET = 13'h0f0c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_88_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_88_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_88_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_89_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_89_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_89_BYTE_OFFSET = 13'h0f10;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_89_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_89_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_89_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_90_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_90_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_90_BYTE_OFFSET = 13'h0f14;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_90_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_90_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_90_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_91_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_91_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_91_BYTE_OFFSET = 13'h0f18;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_91_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_91_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_91_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_92_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_92_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_92_BYTE_OFFSET = 13'h0f1c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_92_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_92_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_92_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_93_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_93_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_93_BYTE_OFFSET = 13'h0f20;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_93_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_93_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_93_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_94_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_94_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_94_BYTE_OFFSET = 13'h0f24;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_94_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_94_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_94_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_95_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_95_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_95_BYTE_OFFSET = 13'h0f28;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_95_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_95_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_95_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_96_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_96_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_96_BYTE_OFFSET = 13'h0f2c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_96_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_96_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_96_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_97_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_97_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_97_BYTE_OFFSET = 13'h0f30;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_97_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_97_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_97_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_98_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_98_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_98_BYTE_OFFSET = 13'h0f34;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_98_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_98_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_98_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_99_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_99_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_99_BYTE_OFFSET = 13'h0f38;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_99_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_99_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_99_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_100_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_100_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_100_BYTE_OFFSET = 13'h0f3c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_100_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_100_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_100_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_101_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_101_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_101_BYTE_OFFSET = 13'h0f40;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_101_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_101_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_101_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_102_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_102_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_102_BYTE_OFFSET = 13'h0f44;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_102_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_102_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_102_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_103_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_103_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_103_BYTE_OFFSET = 13'h0f48;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_103_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_103_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_103_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_104_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_104_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_104_BYTE_OFFSET = 13'h0f4c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_104_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_104_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_104_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_105_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_105_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_105_BYTE_OFFSET = 13'h0f50;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_105_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_105_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_105_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_106_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_106_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_106_BYTE_OFFSET = 13'h0f54;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_106_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_106_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_106_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_107_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_107_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_107_BYTE_OFFSET = 13'h0f58;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_107_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_107_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_107_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_108_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_108_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_108_BYTE_OFFSET = 13'h0f5c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_108_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_108_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_108_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_109_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_109_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_109_BYTE_OFFSET = 13'h0f60;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_109_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_109_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_109_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_110_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_110_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_110_BYTE_OFFSET = 13'h0f64;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_110_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_110_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_110_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_111_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_111_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_111_BYTE_OFFSET = 13'h0f68;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_111_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_111_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_111_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_112_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_112_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_112_BYTE_OFFSET = 13'h0f6c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_112_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_112_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_112_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_113_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_113_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_113_BYTE_OFFSET = 13'h0f70;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_113_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_113_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_113_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_114_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_114_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_114_BYTE_OFFSET = 13'h0f74;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_114_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_114_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_114_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_115_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_115_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_115_BYTE_OFFSET = 13'h0f78;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_115_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_115_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_115_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_116_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_116_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_116_BYTE_OFFSET = 13'h0f7c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_116_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_116_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_116_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_117_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_117_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_117_BYTE_OFFSET = 13'h0f80;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_117_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_117_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_117_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_118_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_118_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_118_BYTE_OFFSET = 13'h0f84;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_118_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_118_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_118_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_119_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_119_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_119_BYTE_OFFSET = 13'h0f88;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_119_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_119_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_119_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_120_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_120_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_120_BYTE_OFFSET = 13'h0f8c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_120_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_120_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_120_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_121_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_121_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_121_BYTE_OFFSET = 13'h0f90;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_121_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_121_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_121_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_122_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_122_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_122_BYTE_OFFSET = 13'h0f94;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_122_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_122_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_122_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_123_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_123_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_123_BYTE_OFFSET = 13'h0f98;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_123_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_123_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_123_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_124_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_124_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_124_BYTE_OFFSET = 13'h0f9c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_124_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_124_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_124_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_125_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_125_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_125_BYTE_OFFSET = 13'h0fa0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_125_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_125_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_125_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_126_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_126_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_126_BYTE_OFFSET = 13'h0fa4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_126_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_126_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_126_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_127_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_127_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_127_BYTE_OFFSET = 13'h0fa8;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_127_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_127_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_127_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_128_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_128_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_128_BYTE_OFFSET = 13'h0fac;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_128_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_128_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_128_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_129_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_129_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_129_BYTE_OFFSET = 13'h0fb0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_129_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_129_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_129_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_130_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_130_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_130_BYTE_OFFSET = 13'h0fb4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_130_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_130_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_130_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_131_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_131_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_131_BYTE_OFFSET = 13'h0fb8;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_131_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_131_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_131_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_132_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_132_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_132_BYTE_OFFSET = 13'h0fbc;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_132_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_132_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_132_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_133_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_133_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_133_BYTE_OFFSET = 13'h0fc0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_133_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_133_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_133_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_134_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_134_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_134_BYTE_OFFSET = 13'h0fc4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_134_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_134_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_134_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_135_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_135_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_135_BYTE_OFFSET = 13'h0fc8;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_135_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_135_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_135_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_136_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_136_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_136_BYTE_OFFSET = 13'h0fcc;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_136_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_136_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_136_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_137_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_137_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_137_BYTE_OFFSET = 13'h0fd0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_137_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_137_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_137_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_138_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_138_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_138_BYTE_OFFSET = 13'h0fd4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_138_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_138_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_138_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_139_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_139_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_139_BYTE_OFFSET = 13'h0fd8;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_139_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_139_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_139_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_140_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_140_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_140_BYTE_OFFSET = 13'h0fdc;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_140_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_140_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_140_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_141_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_141_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_141_BYTE_OFFSET = 13'h0fe0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_141_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_141_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_141_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_142_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_142_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_142_BYTE_OFFSET = 13'h0fe4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_142_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_142_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_142_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_143_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_143_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_143_BYTE_OFFSET = 13'h0fe8;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_143_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_143_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_143_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_144_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_144_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_144_BYTE_OFFSET = 13'h0fec;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_144_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_144_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_144_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_145_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_145_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_145_BYTE_OFFSET = 13'h0ff0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_145_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_145_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_145_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_146_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_146_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_146_BYTE_OFFSET = 13'h0ff4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_146_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_146_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_146_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_147_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_147_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_147_BYTE_OFFSET = 13'h0ff8;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_147_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_147_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_147_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_148_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_148_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_148_BYTE_OFFSET = 13'h0ffc;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_148_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_148_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_148_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_149_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_149_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_149_BYTE_OFFSET = 13'h1000;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_149_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_149_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_149_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_150_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_150_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_150_BYTE_OFFSET = 13'h1004;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_150_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_150_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_150_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_151_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_151_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_151_BYTE_OFFSET = 13'h1008;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_151_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_151_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_151_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_152_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_152_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_152_BYTE_OFFSET = 13'h100c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_152_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_152_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_152_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_153_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_153_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_153_BYTE_OFFSET = 13'h1010;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_153_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_153_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_153_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_154_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_154_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_154_BYTE_OFFSET = 13'h1014;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_154_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_154_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_154_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_155_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_155_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_155_BYTE_OFFSET = 13'h1018;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_155_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_155_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_155_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_156_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_156_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_156_BYTE_OFFSET = 13'h101c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_156_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_156_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_156_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_157_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_157_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_157_BYTE_OFFSET = 13'h1020;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_157_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_157_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_157_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_158_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_158_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_158_BYTE_OFFSET = 13'h1024;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_158_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_158_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_158_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_159_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_159_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_159_BYTE_OFFSET = 13'h1028;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_159_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_159_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_159_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_160_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_160_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_160_BYTE_OFFSET = 13'h102c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_160_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_160_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_160_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_161_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_161_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_161_BYTE_OFFSET = 13'h1030;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_161_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_161_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_161_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_162_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_162_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_162_BYTE_OFFSET = 13'h1034;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_162_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_162_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_162_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_163_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_163_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_163_BYTE_OFFSET = 13'h1038;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_163_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_163_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_163_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_164_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_164_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_164_BYTE_OFFSET = 13'h103c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_164_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_164_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_164_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_165_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_165_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_165_BYTE_OFFSET = 13'h1040;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_165_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_165_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_165_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_166_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_166_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_166_BYTE_OFFSET = 13'h1044;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_166_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_166_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_166_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_167_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_167_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_167_BYTE_OFFSET = 13'h1048;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_167_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_167_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_167_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_168_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_168_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_168_BYTE_OFFSET = 13'h104c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_168_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_168_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_168_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_169_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_169_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_169_BYTE_OFFSET = 13'h1050;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_169_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_169_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_169_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_170_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_170_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_170_BYTE_OFFSET = 13'h1054;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_170_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_170_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_170_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_171_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_171_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_171_BYTE_OFFSET = 13'h1058;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_171_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_171_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_171_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_172_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_172_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_172_BYTE_OFFSET = 13'h105c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_172_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_172_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_172_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_173_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_173_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_173_BYTE_OFFSET = 13'h1060;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_173_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_173_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_173_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_174_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_174_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_174_BYTE_OFFSET = 13'h1064;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_174_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_174_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_174_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_175_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_175_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_175_BYTE_OFFSET = 13'h1068;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_175_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_175_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_175_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_176_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_176_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_176_BYTE_OFFSET = 13'h106c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_176_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_176_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_176_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_177_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_177_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_177_BYTE_OFFSET = 13'h1070;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_177_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_177_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_177_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_178_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_178_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_178_BYTE_OFFSET = 13'h1074;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_178_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_178_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_178_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_179_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_179_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_179_BYTE_OFFSET = 13'h1078;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_179_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_179_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_179_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_180_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_180_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_180_BYTE_OFFSET = 13'h107c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_180_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_180_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_180_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_181_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_181_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_181_BYTE_OFFSET = 13'h1080;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_181_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_181_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_181_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_182_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_182_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_182_BYTE_OFFSET = 13'h1084;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_182_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_182_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_182_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_183_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_183_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_183_BYTE_OFFSET = 13'h1088;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_183_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_183_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_183_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_184_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_184_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_184_BYTE_OFFSET = 13'h108c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_184_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_184_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_184_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_185_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_185_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_185_BYTE_OFFSET = 13'h1090;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_185_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_185_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_185_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_186_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_186_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_186_BYTE_OFFSET = 13'h1094;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_186_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_186_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_186_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_187_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_187_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_187_BYTE_OFFSET = 13'h1098;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_187_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_187_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_187_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_188_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_188_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_188_BYTE_OFFSET = 13'h109c;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_188_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_188_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_188_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_189_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_189_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_189_BYTE_OFFSET = 13'h10a0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_189_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_189_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_189_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_190_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_190_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_190_BYTE_OFFSET = 13'h10a4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_190_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_190_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_190_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_191_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_191_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_191_BYTE_OFFSET = 13'h10a8;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_191_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_191_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_191_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_192_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_192_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_192_BYTE_OFFSET = 13'h10ac;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_192_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_192_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_192_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_193_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_193_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_193_BYTE_OFFSET = 13'h10b0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_193_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_193_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_193_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_194_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_194_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_194_BYTE_OFFSET = 13'h10b4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_194_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_194_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_194_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_195_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_195_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_195_BYTE_OFFSET = 13'h10b8;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_195_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_195_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_195_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_196_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_196_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_196_BYTE_OFFSET = 13'h10bc;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_196_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_196_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_196_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_197_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_197_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_197_BYTE_OFFSET = 13'h10c0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_197_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_197_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_197_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_198_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_198_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_198_BYTE_OFFSET = 13'h10c4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_198_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_198_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_198_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_199_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_199_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_199_BYTE_OFFSET = 13'h10c8;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_199_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_199_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_199_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_200_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_200_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_200_BYTE_OFFSET = 13'h10cc;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_200_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_200_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_200_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_201_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_201_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_201_BYTE_OFFSET = 13'h10d0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_201_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_201_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_201_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_202_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_202_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_202_BYTE_OFFSET = 13'h10d4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_202_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_202_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_202_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_203_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_203_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_203_BYTE_OFFSET = 13'h10d8;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_203_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_203_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_203_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_204_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_204_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_204_BYTE_OFFSET = 13'h10dc;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_204_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_204_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_204_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_205_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_205_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_205_BYTE_OFFSET = 13'h10e0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_205_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_205_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_205_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_206_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_206_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_206_BYTE_OFFSET = 13'h10e4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_206_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_206_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_206_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_207_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_207_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_IN_Q0_1_207_BYTE_OFFSET = 13'h10e8;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_207_CWORD_Q0_1_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_IN_Q0_1_207_CWORD_Q0_1_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_IN_Q0_1_207_CWORD_Q0_1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_ERR_INTRO_DECODER_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_ERR_INTRO_DECODER_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_ERR_INTRO_DECODER_BYTE_OFFSET = 13'h10ec;
  localparam int LDPC_DEC_ERR_INTRO_DECODER_ERR_INTRO_DECODER_BIT_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_ERR_INTRO_DECODER_ERR_INTRO_DECODER_BIT_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_ERR_INTRO_DECODER_ERR_INTRO_DECODER_BIT_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_0_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_0_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_0_BYTE_OFFSET = 13'h10f0;
  localparam int LDPC_DEC_EXPSYND_0_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_0_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_0_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_1_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_1_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_1_BYTE_OFFSET = 13'h10f4;
  localparam int LDPC_DEC_EXPSYND_1_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_1_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_1_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_2_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_2_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_2_BYTE_OFFSET = 13'h10f8;
  localparam int LDPC_DEC_EXPSYND_2_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_2_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_2_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_3_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_3_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_3_BYTE_OFFSET = 13'h10fc;
  localparam int LDPC_DEC_EXPSYND_3_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_3_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_3_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_4_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_4_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_4_BYTE_OFFSET = 13'h1100;
  localparam int LDPC_DEC_EXPSYND_4_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_4_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_4_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_5_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_5_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_5_BYTE_OFFSET = 13'h1104;
  localparam int LDPC_DEC_EXPSYND_5_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_5_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_5_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_6_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_6_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_6_BYTE_OFFSET = 13'h1108;
  localparam int LDPC_DEC_EXPSYND_6_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_6_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_6_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_7_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_7_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_7_BYTE_OFFSET = 13'h110c;
  localparam int LDPC_DEC_EXPSYND_7_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_7_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_7_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_8_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_8_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_8_BYTE_OFFSET = 13'h1110;
  localparam int LDPC_DEC_EXPSYND_8_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_8_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_8_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_9_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_9_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_9_BYTE_OFFSET = 13'h1114;
  localparam int LDPC_DEC_EXPSYND_9_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_9_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_9_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_10_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_10_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_10_BYTE_OFFSET = 13'h1118;
  localparam int LDPC_DEC_EXPSYND_10_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_10_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_10_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_11_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_11_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_11_BYTE_OFFSET = 13'h111c;
  localparam int LDPC_DEC_EXPSYND_11_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_11_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_11_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_12_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_12_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_12_BYTE_OFFSET = 13'h1120;
  localparam int LDPC_DEC_EXPSYND_12_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_12_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_12_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_13_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_13_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_13_BYTE_OFFSET = 13'h1124;
  localparam int LDPC_DEC_EXPSYND_13_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_13_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_13_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_14_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_14_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_14_BYTE_OFFSET = 13'h1128;
  localparam int LDPC_DEC_EXPSYND_14_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_14_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_14_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_15_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_15_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_15_BYTE_OFFSET = 13'h112c;
  localparam int LDPC_DEC_EXPSYND_15_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_15_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_15_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_16_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_16_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_16_BYTE_OFFSET = 13'h1130;
  localparam int LDPC_DEC_EXPSYND_16_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_16_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_16_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_17_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_17_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_17_BYTE_OFFSET = 13'h1134;
  localparam int LDPC_DEC_EXPSYND_17_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_17_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_17_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_18_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_18_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_18_BYTE_OFFSET = 13'h1138;
  localparam int LDPC_DEC_EXPSYND_18_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_18_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_18_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_19_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_19_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_19_BYTE_OFFSET = 13'h113c;
  localparam int LDPC_DEC_EXPSYND_19_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_19_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_19_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_20_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_20_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_20_BYTE_OFFSET = 13'h1140;
  localparam int LDPC_DEC_EXPSYND_20_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_20_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_20_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_21_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_21_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_21_BYTE_OFFSET = 13'h1144;
  localparam int LDPC_DEC_EXPSYND_21_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_21_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_21_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_22_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_22_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_22_BYTE_OFFSET = 13'h1148;
  localparam int LDPC_DEC_EXPSYND_22_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_22_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_22_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_23_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_23_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_23_BYTE_OFFSET = 13'h114c;
  localparam int LDPC_DEC_EXPSYND_23_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_23_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_23_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_24_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_24_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_24_BYTE_OFFSET = 13'h1150;
  localparam int LDPC_DEC_EXPSYND_24_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_24_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_24_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_25_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_25_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_25_BYTE_OFFSET = 13'h1154;
  localparam int LDPC_DEC_EXPSYND_25_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_25_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_25_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_26_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_26_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_26_BYTE_OFFSET = 13'h1158;
  localparam int LDPC_DEC_EXPSYND_26_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_26_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_26_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_27_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_27_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_27_BYTE_OFFSET = 13'h115c;
  localparam int LDPC_DEC_EXPSYND_27_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_27_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_27_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_28_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_28_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_28_BYTE_OFFSET = 13'h1160;
  localparam int LDPC_DEC_EXPSYND_28_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_28_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_28_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_29_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_29_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_29_BYTE_OFFSET = 13'h1164;
  localparam int LDPC_DEC_EXPSYND_29_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_29_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_29_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_30_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_30_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_30_BYTE_OFFSET = 13'h1168;
  localparam int LDPC_DEC_EXPSYND_30_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_30_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_30_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_31_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_31_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_31_BYTE_OFFSET = 13'h116c;
  localparam int LDPC_DEC_EXPSYND_31_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_31_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_31_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_32_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_32_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_32_BYTE_OFFSET = 13'h1170;
  localparam int LDPC_DEC_EXPSYND_32_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_32_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_32_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_33_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_33_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_33_BYTE_OFFSET = 13'h1174;
  localparam int LDPC_DEC_EXPSYND_33_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_33_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_33_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_34_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_34_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_34_BYTE_OFFSET = 13'h1178;
  localparam int LDPC_DEC_EXPSYND_34_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_34_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_34_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_35_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_35_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_35_BYTE_OFFSET = 13'h117c;
  localparam int LDPC_DEC_EXPSYND_35_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_35_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_35_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_36_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_36_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_36_BYTE_OFFSET = 13'h1180;
  localparam int LDPC_DEC_EXPSYND_36_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_36_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_36_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_37_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_37_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_37_BYTE_OFFSET = 13'h1184;
  localparam int LDPC_DEC_EXPSYND_37_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_37_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_37_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_38_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_38_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_38_BYTE_OFFSET = 13'h1188;
  localparam int LDPC_DEC_EXPSYND_38_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_38_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_38_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_39_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_39_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_39_BYTE_OFFSET = 13'h118c;
  localparam int LDPC_DEC_EXPSYND_39_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_39_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_39_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_40_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_40_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_40_BYTE_OFFSET = 13'h1190;
  localparam int LDPC_DEC_EXPSYND_40_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_40_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_40_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_41_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_41_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_41_BYTE_OFFSET = 13'h1194;
  localparam int LDPC_DEC_EXPSYND_41_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_41_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_41_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_42_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_42_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_42_BYTE_OFFSET = 13'h1198;
  localparam int LDPC_DEC_EXPSYND_42_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_42_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_42_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_43_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_43_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_43_BYTE_OFFSET = 13'h119c;
  localparam int LDPC_DEC_EXPSYND_43_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_43_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_43_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_44_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_44_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_44_BYTE_OFFSET = 13'h11a0;
  localparam int LDPC_DEC_EXPSYND_44_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_44_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_44_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_45_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_45_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_45_BYTE_OFFSET = 13'h11a4;
  localparam int LDPC_DEC_EXPSYND_45_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_45_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_45_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_46_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_46_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_46_BYTE_OFFSET = 13'h11a8;
  localparam int LDPC_DEC_EXPSYND_46_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_46_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_46_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_47_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_47_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_47_BYTE_OFFSET = 13'h11ac;
  localparam int LDPC_DEC_EXPSYND_47_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_47_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_47_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_48_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_48_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_48_BYTE_OFFSET = 13'h11b0;
  localparam int LDPC_DEC_EXPSYND_48_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_48_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_48_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_49_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_49_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_49_BYTE_OFFSET = 13'h11b4;
  localparam int LDPC_DEC_EXPSYND_49_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_49_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_49_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_50_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_50_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_50_BYTE_OFFSET = 13'h11b8;
  localparam int LDPC_DEC_EXPSYND_50_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_50_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_50_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_51_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_51_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_51_BYTE_OFFSET = 13'h11bc;
  localparam int LDPC_DEC_EXPSYND_51_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_51_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_51_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_52_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_52_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_52_BYTE_OFFSET = 13'h11c0;
  localparam int LDPC_DEC_EXPSYND_52_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_52_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_52_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_53_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_53_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_53_BYTE_OFFSET = 13'h11c4;
  localparam int LDPC_DEC_EXPSYND_53_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_53_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_53_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_54_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_54_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_54_BYTE_OFFSET = 13'h11c8;
  localparam int LDPC_DEC_EXPSYND_54_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_54_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_54_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_55_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_55_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_55_BYTE_OFFSET = 13'h11cc;
  localparam int LDPC_DEC_EXPSYND_55_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_55_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_55_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_56_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_56_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_56_BYTE_OFFSET = 13'h11d0;
  localparam int LDPC_DEC_EXPSYND_56_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_56_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_56_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_57_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_57_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_57_BYTE_OFFSET = 13'h11d4;
  localparam int LDPC_DEC_EXPSYND_57_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_57_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_57_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_58_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_58_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_58_BYTE_OFFSET = 13'h11d8;
  localparam int LDPC_DEC_EXPSYND_58_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_58_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_58_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_59_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_59_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_59_BYTE_OFFSET = 13'h11dc;
  localparam int LDPC_DEC_EXPSYND_59_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_59_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_59_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_60_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_60_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_60_BYTE_OFFSET = 13'h11e0;
  localparam int LDPC_DEC_EXPSYND_60_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_60_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_60_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_61_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_61_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_61_BYTE_OFFSET = 13'h11e4;
  localparam int LDPC_DEC_EXPSYND_61_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_61_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_61_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_62_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_62_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_62_BYTE_OFFSET = 13'h11e8;
  localparam int LDPC_DEC_EXPSYND_62_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_62_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_62_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_63_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_63_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_63_BYTE_OFFSET = 13'h11ec;
  localparam int LDPC_DEC_EXPSYND_63_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_63_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_63_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_64_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_64_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_64_BYTE_OFFSET = 13'h11f0;
  localparam int LDPC_DEC_EXPSYND_64_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_64_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_64_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_65_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_65_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_65_BYTE_OFFSET = 13'h11f4;
  localparam int LDPC_DEC_EXPSYND_65_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_65_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_65_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_66_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_66_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_66_BYTE_OFFSET = 13'h11f8;
  localparam int LDPC_DEC_EXPSYND_66_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_66_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_66_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_67_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_67_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_67_BYTE_OFFSET = 13'h11fc;
  localparam int LDPC_DEC_EXPSYND_67_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_67_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_67_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_68_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_68_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_68_BYTE_OFFSET = 13'h1200;
  localparam int LDPC_DEC_EXPSYND_68_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_68_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_68_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_69_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_69_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_69_BYTE_OFFSET = 13'h1204;
  localparam int LDPC_DEC_EXPSYND_69_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_69_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_69_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_70_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_70_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_70_BYTE_OFFSET = 13'h1208;
  localparam int LDPC_DEC_EXPSYND_70_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_70_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_70_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_71_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_71_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_71_BYTE_OFFSET = 13'h120c;
  localparam int LDPC_DEC_EXPSYND_71_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_71_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_71_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_72_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_72_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_72_BYTE_OFFSET = 13'h1210;
  localparam int LDPC_DEC_EXPSYND_72_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_72_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_72_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_73_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_73_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_73_BYTE_OFFSET = 13'h1214;
  localparam int LDPC_DEC_EXPSYND_73_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_73_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_73_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_74_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_74_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_74_BYTE_OFFSET = 13'h1218;
  localparam int LDPC_DEC_EXPSYND_74_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_74_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_74_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_75_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_75_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_75_BYTE_OFFSET = 13'h121c;
  localparam int LDPC_DEC_EXPSYND_75_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_75_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_75_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_76_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_76_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_76_BYTE_OFFSET = 13'h1220;
  localparam int LDPC_DEC_EXPSYND_76_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_76_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_76_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_77_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_77_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_77_BYTE_OFFSET = 13'h1224;
  localparam int LDPC_DEC_EXPSYND_77_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_77_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_77_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_78_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_78_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_78_BYTE_OFFSET = 13'h1228;
  localparam int LDPC_DEC_EXPSYND_78_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_78_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_78_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_79_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_79_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_79_BYTE_OFFSET = 13'h122c;
  localparam int LDPC_DEC_EXPSYND_79_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_79_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_79_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_80_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_80_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_80_BYTE_OFFSET = 13'h1230;
  localparam int LDPC_DEC_EXPSYND_80_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_80_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_80_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_81_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_81_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_81_BYTE_OFFSET = 13'h1234;
  localparam int LDPC_DEC_EXPSYND_81_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_81_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_81_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_82_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_82_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_82_BYTE_OFFSET = 13'h1238;
  localparam int LDPC_DEC_EXPSYND_82_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_82_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_82_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_83_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_83_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_83_BYTE_OFFSET = 13'h123c;
  localparam int LDPC_DEC_EXPSYND_83_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_83_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_83_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_84_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_84_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_84_BYTE_OFFSET = 13'h1240;
  localparam int LDPC_DEC_EXPSYND_84_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_84_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_84_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_85_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_85_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_85_BYTE_OFFSET = 13'h1244;
  localparam int LDPC_DEC_EXPSYND_85_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_85_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_85_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_86_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_86_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_86_BYTE_OFFSET = 13'h1248;
  localparam int LDPC_DEC_EXPSYND_86_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_86_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_86_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_87_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_87_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_87_BYTE_OFFSET = 13'h124c;
  localparam int LDPC_DEC_EXPSYND_87_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_87_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_87_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_88_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_88_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_88_BYTE_OFFSET = 13'h1250;
  localparam int LDPC_DEC_EXPSYND_88_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_88_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_88_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_89_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_89_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_89_BYTE_OFFSET = 13'h1254;
  localparam int LDPC_DEC_EXPSYND_89_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_89_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_89_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_90_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_90_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_90_BYTE_OFFSET = 13'h1258;
  localparam int LDPC_DEC_EXPSYND_90_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_90_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_90_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_91_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_91_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_91_BYTE_OFFSET = 13'h125c;
  localparam int LDPC_DEC_EXPSYND_91_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_91_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_91_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_92_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_92_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_92_BYTE_OFFSET = 13'h1260;
  localparam int LDPC_DEC_EXPSYND_92_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_92_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_92_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_93_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_93_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_93_BYTE_OFFSET = 13'h1264;
  localparam int LDPC_DEC_EXPSYND_93_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_93_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_93_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_94_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_94_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_94_BYTE_OFFSET = 13'h1268;
  localparam int LDPC_DEC_EXPSYND_94_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_94_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_94_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_95_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_95_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_95_BYTE_OFFSET = 13'h126c;
  localparam int LDPC_DEC_EXPSYND_95_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_95_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_95_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_96_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_96_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_96_BYTE_OFFSET = 13'h1270;
  localparam int LDPC_DEC_EXPSYND_96_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_96_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_96_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_97_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_97_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_97_BYTE_OFFSET = 13'h1274;
  localparam int LDPC_DEC_EXPSYND_97_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_97_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_97_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_98_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_98_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_98_BYTE_OFFSET = 13'h1278;
  localparam int LDPC_DEC_EXPSYND_98_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_98_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_98_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_99_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_99_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_99_BYTE_OFFSET = 13'h127c;
  localparam int LDPC_DEC_EXPSYND_99_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_99_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_99_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_100_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_100_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_100_BYTE_OFFSET = 13'h1280;
  localparam int LDPC_DEC_EXPSYND_100_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_100_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_100_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_101_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_101_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_101_BYTE_OFFSET = 13'h1284;
  localparam int LDPC_DEC_EXPSYND_101_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_101_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_101_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_102_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_102_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_102_BYTE_OFFSET = 13'h1288;
  localparam int LDPC_DEC_EXPSYND_102_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_102_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_102_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_103_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_103_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_103_BYTE_OFFSET = 13'h128c;
  localparam int LDPC_DEC_EXPSYND_103_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_103_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_103_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_104_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_104_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_104_BYTE_OFFSET = 13'h1290;
  localparam int LDPC_DEC_EXPSYND_104_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_104_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_104_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_105_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_105_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_105_BYTE_OFFSET = 13'h1294;
  localparam int LDPC_DEC_EXPSYND_105_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_105_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_105_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_106_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_106_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_106_BYTE_OFFSET = 13'h1298;
  localparam int LDPC_DEC_EXPSYND_106_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_106_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_106_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_107_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_107_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_107_BYTE_OFFSET = 13'h129c;
  localparam int LDPC_DEC_EXPSYND_107_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_107_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_107_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_108_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_108_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_108_BYTE_OFFSET = 13'h12a0;
  localparam int LDPC_DEC_EXPSYND_108_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_108_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_108_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_109_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_109_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_109_BYTE_OFFSET = 13'h12a4;
  localparam int LDPC_DEC_EXPSYND_109_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_109_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_109_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_110_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_110_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_110_BYTE_OFFSET = 13'h12a8;
  localparam int LDPC_DEC_EXPSYND_110_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_110_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_110_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_111_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_111_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_111_BYTE_OFFSET = 13'h12ac;
  localparam int LDPC_DEC_EXPSYND_111_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_111_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_111_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_112_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_112_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_112_BYTE_OFFSET = 13'h12b0;
  localparam int LDPC_DEC_EXPSYND_112_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_112_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_112_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_113_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_113_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_113_BYTE_OFFSET = 13'h12b4;
  localparam int LDPC_DEC_EXPSYND_113_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_113_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_113_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_114_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_114_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_114_BYTE_OFFSET = 13'h12b8;
  localparam int LDPC_DEC_EXPSYND_114_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_114_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_114_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_115_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_115_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_115_BYTE_OFFSET = 13'h12bc;
  localparam int LDPC_DEC_EXPSYND_115_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_115_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_115_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_116_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_116_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_116_BYTE_OFFSET = 13'h12c0;
  localparam int LDPC_DEC_EXPSYND_116_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_116_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_116_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_117_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_117_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_117_BYTE_OFFSET = 13'h12c4;
  localparam int LDPC_DEC_EXPSYND_117_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_117_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_117_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_118_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_118_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_118_BYTE_OFFSET = 13'h12c8;
  localparam int LDPC_DEC_EXPSYND_118_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_118_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_118_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_119_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_119_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_119_BYTE_OFFSET = 13'h12cc;
  localparam int LDPC_DEC_EXPSYND_119_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_119_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_119_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_120_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_120_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_120_BYTE_OFFSET = 13'h12d0;
  localparam int LDPC_DEC_EXPSYND_120_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_120_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_120_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_121_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_121_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_121_BYTE_OFFSET = 13'h12d4;
  localparam int LDPC_DEC_EXPSYND_121_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_121_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_121_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_122_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_122_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_122_BYTE_OFFSET = 13'h12d8;
  localparam int LDPC_DEC_EXPSYND_122_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_122_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_122_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_123_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_123_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_123_BYTE_OFFSET = 13'h12dc;
  localparam int LDPC_DEC_EXPSYND_123_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_123_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_123_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_124_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_124_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_124_BYTE_OFFSET = 13'h12e0;
  localparam int LDPC_DEC_EXPSYND_124_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_124_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_124_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_125_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_125_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_125_BYTE_OFFSET = 13'h12e4;
  localparam int LDPC_DEC_EXPSYND_125_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_125_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_125_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_126_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_126_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_126_BYTE_OFFSET = 13'h12e8;
  localparam int LDPC_DEC_EXPSYND_126_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_126_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_126_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_127_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_127_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_127_BYTE_OFFSET = 13'h12ec;
  localparam int LDPC_DEC_EXPSYND_127_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_127_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_127_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_128_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_128_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_128_BYTE_OFFSET = 13'h12f0;
  localparam int LDPC_DEC_EXPSYND_128_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_128_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_128_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_129_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_129_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_129_BYTE_OFFSET = 13'h12f4;
  localparam int LDPC_DEC_EXPSYND_129_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_129_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_129_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_130_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_130_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_130_BYTE_OFFSET = 13'h12f8;
  localparam int LDPC_DEC_EXPSYND_130_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_130_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_130_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_131_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_131_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_131_BYTE_OFFSET = 13'h12fc;
  localparam int LDPC_DEC_EXPSYND_131_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_131_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_131_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_132_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_132_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_132_BYTE_OFFSET = 13'h1300;
  localparam int LDPC_DEC_EXPSYND_132_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_132_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_132_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_133_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_133_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_133_BYTE_OFFSET = 13'h1304;
  localparam int LDPC_DEC_EXPSYND_133_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_133_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_133_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_134_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_134_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_134_BYTE_OFFSET = 13'h1308;
  localparam int LDPC_DEC_EXPSYND_134_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_134_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_134_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_135_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_135_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_135_BYTE_OFFSET = 13'h130c;
  localparam int LDPC_DEC_EXPSYND_135_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_135_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_135_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_136_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_136_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_136_BYTE_OFFSET = 13'h1310;
  localparam int LDPC_DEC_EXPSYND_136_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_136_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_136_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_137_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_137_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_137_BYTE_OFFSET = 13'h1314;
  localparam int LDPC_DEC_EXPSYND_137_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_137_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_137_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_138_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_138_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_138_BYTE_OFFSET = 13'h1318;
  localparam int LDPC_DEC_EXPSYND_138_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_138_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_138_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_139_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_139_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_139_BYTE_OFFSET = 13'h131c;
  localparam int LDPC_DEC_EXPSYND_139_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_139_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_139_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_140_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_140_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_140_BYTE_OFFSET = 13'h1320;
  localparam int LDPC_DEC_EXPSYND_140_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_140_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_140_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_141_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_141_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_141_BYTE_OFFSET = 13'h1324;
  localparam int LDPC_DEC_EXPSYND_141_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_141_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_141_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_142_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_142_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_142_BYTE_OFFSET = 13'h1328;
  localparam int LDPC_DEC_EXPSYND_142_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_142_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_142_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_143_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_143_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_143_BYTE_OFFSET = 13'h132c;
  localparam int LDPC_DEC_EXPSYND_143_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_143_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_143_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_144_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_144_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_144_BYTE_OFFSET = 13'h1330;
  localparam int LDPC_DEC_EXPSYND_144_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_144_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_144_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_145_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_145_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_145_BYTE_OFFSET = 13'h1334;
  localparam int LDPC_DEC_EXPSYND_145_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_145_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_145_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_146_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_146_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_146_BYTE_OFFSET = 13'h1338;
  localparam int LDPC_DEC_EXPSYND_146_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_146_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_146_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_147_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_147_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_147_BYTE_OFFSET = 13'h133c;
  localparam int LDPC_DEC_EXPSYND_147_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_147_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_147_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_148_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_148_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_148_BYTE_OFFSET = 13'h1340;
  localparam int LDPC_DEC_EXPSYND_148_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_148_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_148_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_149_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_149_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_149_BYTE_OFFSET = 13'h1344;
  localparam int LDPC_DEC_EXPSYND_149_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_149_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_149_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_150_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_150_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_150_BYTE_OFFSET = 13'h1348;
  localparam int LDPC_DEC_EXPSYND_150_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_150_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_150_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_151_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_151_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_151_BYTE_OFFSET = 13'h134c;
  localparam int LDPC_DEC_EXPSYND_151_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_151_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_151_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_152_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_152_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_152_BYTE_OFFSET = 13'h1350;
  localparam int LDPC_DEC_EXPSYND_152_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_152_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_152_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_153_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_153_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_153_BYTE_OFFSET = 13'h1354;
  localparam int LDPC_DEC_EXPSYND_153_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_153_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_153_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_154_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_154_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_154_BYTE_OFFSET = 13'h1358;
  localparam int LDPC_DEC_EXPSYND_154_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_154_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_154_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_155_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_155_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_155_BYTE_OFFSET = 13'h135c;
  localparam int LDPC_DEC_EXPSYND_155_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_155_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_155_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_156_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_156_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_156_BYTE_OFFSET = 13'h1360;
  localparam int LDPC_DEC_EXPSYND_156_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_156_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_156_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_157_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_157_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_157_BYTE_OFFSET = 13'h1364;
  localparam int LDPC_DEC_EXPSYND_157_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_157_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_157_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_158_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_158_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_158_BYTE_OFFSET = 13'h1368;
  localparam int LDPC_DEC_EXPSYND_158_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_158_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_158_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_159_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_159_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_159_BYTE_OFFSET = 13'h136c;
  localparam int LDPC_DEC_EXPSYND_159_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_159_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_159_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_160_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_160_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_160_BYTE_OFFSET = 13'h1370;
  localparam int LDPC_DEC_EXPSYND_160_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_160_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_160_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_161_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_161_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_161_BYTE_OFFSET = 13'h1374;
  localparam int LDPC_DEC_EXPSYND_161_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_161_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_161_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_162_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_162_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_162_BYTE_OFFSET = 13'h1378;
  localparam int LDPC_DEC_EXPSYND_162_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_162_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_162_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_163_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_163_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_163_BYTE_OFFSET = 13'h137c;
  localparam int LDPC_DEC_EXPSYND_163_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_163_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_163_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_164_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_164_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_164_BYTE_OFFSET = 13'h1380;
  localparam int LDPC_DEC_EXPSYND_164_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_164_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_164_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_165_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_165_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_165_BYTE_OFFSET = 13'h1384;
  localparam int LDPC_DEC_EXPSYND_165_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_165_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_165_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_166_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_166_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_166_BYTE_OFFSET = 13'h1388;
  localparam int LDPC_DEC_EXPSYND_166_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_166_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_166_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_EXPSYND_167_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_EXPSYND_167_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_EXPSYND_167_BYTE_OFFSET = 13'h138c;
  localparam int LDPC_DEC_EXPSYND_167_EXP_SYN_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_EXPSYND_167_EXP_SYN_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_EXPSYND_167_EXP_SYN_BIT_OFFSET = 0;
  localparam int LDPC_DEC_PROBABILITY_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_PROBABILITY_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_PROBABILITY_BYTE_OFFSET = 13'h1390;
  localparam int LDPC_DEC_PROBABILITY_PERC_PROBABILITY_BIT_WIDTH = 32;
  localparam bit [31:0] LDPC_DEC_PROBABILITY_PERC_PROBABILITY_BIT_MASK = 32'hffffffff;
  localparam int LDPC_DEC_PROBABILITY_PERC_PROBABILITY_BIT_OFFSET = 0;
  localparam int LDPC_DEC_HAMDIST_LOOP_MAX_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_HAMDIST_LOOP_MAX_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_HAMDIST_LOOP_MAX_BYTE_OFFSET = 13'h1394;
  localparam int LDPC_DEC_HAMDIST_LOOP_MAX_HAMDIST_LOOP_MAX_BIT_WIDTH = 32;
  localparam bit [31:0] LDPC_DEC_HAMDIST_LOOP_MAX_HAMDIST_LOOP_MAX_BIT_MASK = 32'hffffffff;
  localparam int LDPC_DEC_HAMDIST_LOOP_MAX_HAMDIST_LOOP_MAX_BIT_OFFSET = 0;
  localparam int LDPC_DEC_HAMDIST_LOOP_PERCENTAGE_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_HAMDIST_LOOP_PERCENTAGE_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_HAMDIST_LOOP_PERCENTAGE_BYTE_OFFSET = 13'h1398;
  localparam int LDPC_DEC_HAMDIST_LOOP_PERCENTAGE_HAMDIST_LOOP_PERCENTAGE_BIT_WIDTH = 32;
  localparam bit [31:0] LDPC_DEC_HAMDIST_LOOP_PERCENTAGE_HAMDIST_LOOP_PERCENTAGE_BIT_MASK = 32'hffffffff;
  localparam int LDPC_DEC_HAMDIST_LOOP_PERCENTAGE_HAMDIST_LOOP_PERCENTAGE_BIT_OFFSET = 0;
  localparam int LDPC_DEC_HAMDIST_IIR1_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_HAMDIST_IIR1_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_HAMDIST_IIR1_BYTE_OFFSET = 13'h139c;
  localparam int LDPC_DEC_HAMDIST_IIR1_HAMDIST_IIR1_BIT_WIDTH = 32;
  localparam bit [31:0] LDPC_DEC_HAMDIST_IIR1_HAMDIST_IIR1_BIT_MASK = 32'hffffffff;
  localparam int LDPC_DEC_HAMDIST_IIR1_HAMDIST_IIR1_BIT_OFFSET = 0;
  localparam int LDPC_DEC_HAMDIST_IIR2_NOT_USED_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_HAMDIST_IIR2_NOT_USED_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_HAMDIST_IIR2_NOT_USED_BYTE_OFFSET = 13'h13a0;
  localparam int LDPC_DEC_HAMDIST_IIR2_NOT_USED_HAMDIST_IIR2_BIT_WIDTH = 32;
  localparam bit [31:0] LDPC_DEC_HAMDIST_IIR2_NOT_USED_HAMDIST_IIR2_BIT_MASK = 32'hffffffff;
  localparam int LDPC_DEC_HAMDIST_IIR2_NOT_USED_HAMDIST_IIR2_BIT_OFFSET = 0;
  localparam int LDPC_DEC_HAMDIST_IIR3_NOT_USED_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_HAMDIST_IIR3_NOT_USED_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_HAMDIST_IIR3_NOT_USED_BYTE_OFFSET = 13'h13a4;
  localparam int LDPC_DEC_HAMDIST_IIR3_NOT_USED_HAMDIST_IIR3_BIT_WIDTH = 32;
  localparam bit [31:0] LDPC_DEC_HAMDIST_IIR3_NOT_USED_HAMDIST_IIR3_BIT_MASK = 32'hffffffff;
  localparam int LDPC_DEC_HAMDIST_IIR3_NOT_USED_HAMDIST_IIR3_BIT_OFFSET = 0;
  localparam int LDPC_DEC_SYN_VALID_CWORD_DEC_FINAL_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_SYN_VALID_CWORD_DEC_FINAL_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_SYN_VALID_CWORD_DEC_FINAL_BYTE_OFFSET = 13'h13a8;
  localparam int LDPC_DEC_SYN_VALID_CWORD_DEC_FINAL_SYN_VALID_CWORD_DEC_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_SYN_VALID_CWORD_DEC_FINAL_SYN_VALID_CWORD_DEC_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_SYN_VALID_CWORD_DEC_FINAL_SYN_VALID_CWORD_DEC_BIT_OFFSET = 0;
  localparam int LDPC_DEC_START_DEC_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_START_DEC_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_START_DEC_BYTE_OFFSET = 13'h13ac;
  localparam int LDPC_DEC_START_DEC_START_DEC_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_START_DEC_START_DEC_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_START_DEC_START_DEC_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CONVERGED_LOOPS_ENDED_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CONVERGED_LOOPS_ENDED_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CONVERGED_LOOPS_ENDED_BYTE_OFFSET = 13'h13b0;
  localparam int LDPC_DEC_CONVERGED_LOOPS_ENDED_CONVERGED_LOOPS_ENDED_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CONVERGED_LOOPS_ENDED_CONVERGED_LOOPS_ENDED_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CONVERGED_LOOPS_ENDED_CONVERGED_LOOPS_ENDED_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CONVERGED_PASS_FAIL_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CONVERGED_PASS_FAIL_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CONVERGED_PASS_FAIL_BYTE_OFFSET = 13'h13b4;
  localparam int LDPC_DEC_CONVERGED_PASS_FAIL_CONVERGED_PASS_FAIL_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CONVERGED_PASS_FAIL_CONVERGED_PASS_FAIL_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CONVERGED_PASS_FAIL_CONVERGED_PASS_FAIL_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_0_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_0_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_0_BYTE_OFFSET = 13'h13b8;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_0_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_0_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_0_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_1_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_1_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_1_BYTE_OFFSET = 13'h13bc;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_1_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_1_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_1_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_2_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_2_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_2_BYTE_OFFSET = 13'h13c0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_2_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_2_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_2_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_3_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_3_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_3_BYTE_OFFSET = 13'h13c4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_3_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_3_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_3_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_4_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_4_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_4_BYTE_OFFSET = 13'h13c8;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_4_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_4_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_4_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_5_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_5_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_5_BYTE_OFFSET = 13'h13cc;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_5_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_5_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_5_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_6_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_6_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_6_BYTE_OFFSET = 13'h13d0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_6_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_6_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_6_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_7_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_7_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_7_BYTE_OFFSET = 13'h13d4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_7_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_7_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_7_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_8_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_8_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_8_BYTE_OFFSET = 13'h13d8;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_8_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_8_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_8_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_9_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_9_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_9_BYTE_OFFSET = 13'h13dc;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_9_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_9_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_9_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_10_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_10_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_10_BYTE_OFFSET = 13'h13e0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_10_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_10_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_10_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_11_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_11_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_11_BYTE_OFFSET = 13'h13e4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_11_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_11_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_11_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_12_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_12_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_12_BYTE_OFFSET = 13'h13e8;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_12_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_12_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_12_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_13_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_13_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_13_BYTE_OFFSET = 13'h13ec;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_13_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_13_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_13_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_14_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_14_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_14_BYTE_OFFSET = 13'h13f0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_14_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_14_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_14_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_15_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_15_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_15_BYTE_OFFSET = 13'h13f4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_15_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_15_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_15_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_16_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_16_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_16_BYTE_OFFSET = 13'h13f8;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_16_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_16_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_16_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_17_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_17_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_17_BYTE_OFFSET = 13'h13fc;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_17_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_17_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_17_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_18_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_18_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_18_BYTE_OFFSET = 13'h1400;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_18_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_18_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_18_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_19_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_19_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_19_BYTE_OFFSET = 13'h1404;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_19_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_19_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_19_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_20_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_20_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_20_BYTE_OFFSET = 13'h1408;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_20_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_20_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_20_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_21_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_21_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_21_BYTE_OFFSET = 13'h140c;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_21_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_21_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_21_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_22_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_22_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_22_BYTE_OFFSET = 13'h1410;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_22_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_22_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_22_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_23_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_23_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_23_BYTE_OFFSET = 13'h1414;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_23_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_23_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_23_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_24_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_24_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_24_BYTE_OFFSET = 13'h1418;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_24_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_24_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_24_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_25_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_25_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_25_BYTE_OFFSET = 13'h141c;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_25_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_25_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_25_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_26_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_26_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_26_BYTE_OFFSET = 13'h1420;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_26_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_26_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_26_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_27_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_27_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_27_BYTE_OFFSET = 13'h1424;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_27_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_27_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_27_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_28_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_28_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_28_BYTE_OFFSET = 13'h1428;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_28_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_28_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_28_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_29_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_29_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_29_BYTE_OFFSET = 13'h142c;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_29_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_29_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_29_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_30_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_30_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_30_BYTE_OFFSET = 13'h1430;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_30_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_30_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_30_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_31_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_31_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_31_BYTE_OFFSET = 13'h1434;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_31_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_31_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_31_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_32_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_32_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_32_BYTE_OFFSET = 13'h1438;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_32_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_32_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_32_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_33_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_33_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_33_BYTE_OFFSET = 13'h143c;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_33_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_33_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_33_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_34_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_34_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_34_BYTE_OFFSET = 13'h1440;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_34_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_34_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_34_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_35_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_35_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_35_BYTE_OFFSET = 13'h1444;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_35_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_35_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_35_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_36_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_36_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_36_BYTE_OFFSET = 13'h1448;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_36_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_36_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_36_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_37_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_37_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_37_BYTE_OFFSET = 13'h144c;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_37_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_37_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_37_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_38_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_38_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_38_BYTE_OFFSET = 13'h1450;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_38_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_38_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_38_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_39_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_39_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_39_BYTE_OFFSET = 13'h1454;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_39_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_39_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_39_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_40_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_40_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_40_BYTE_OFFSET = 13'h1458;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_40_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_40_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_40_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_41_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_41_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_41_BYTE_OFFSET = 13'h145c;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_41_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_41_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_41_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_42_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_42_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_42_BYTE_OFFSET = 13'h1460;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_42_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_42_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_42_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_43_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_43_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_43_BYTE_OFFSET = 13'h1464;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_43_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_43_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_43_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_44_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_44_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_44_BYTE_OFFSET = 13'h1468;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_44_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_44_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_44_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_45_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_45_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_45_BYTE_OFFSET = 13'h146c;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_45_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_45_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_45_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_46_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_46_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_46_BYTE_OFFSET = 13'h1470;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_46_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_46_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_46_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_47_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_47_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_47_BYTE_OFFSET = 13'h1474;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_47_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_47_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_47_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_48_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_48_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_48_BYTE_OFFSET = 13'h1478;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_48_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_48_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_48_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_49_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_49_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_49_BYTE_OFFSET = 13'h147c;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_49_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_49_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_49_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_50_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_50_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_50_BYTE_OFFSET = 13'h1480;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_50_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_50_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_50_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_51_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_51_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_51_BYTE_OFFSET = 13'h1484;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_51_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_51_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_51_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_52_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_52_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_52_BYTE_OFFSET = 13'h1488;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_52_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_52_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_52_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_53_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_53_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_53_BYTE_OFFSET = 13'h148c;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_53_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_53_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_53_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_54_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_54_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_54_BYTE_OFFSET = 13'h1490;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_54_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_54_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_54_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_55_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_55_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_55_BYTE_OFFSET = 13'h1494;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_55_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_55_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_55_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_56_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_56_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_56_BYTE_OFFSET = 13'h1498;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_56_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_56_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_56_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_57_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_57_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_57_BYTE_OFFSET = 13'h149c;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_57_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_57_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_57_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_58_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_58_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_58_BYTE_OFFSET = 13'h14a0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_58_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_58_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_58_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_59_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_59_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_59_BYTE_OFFSET = 13'h14a4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_59_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_59_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_59_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_60_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_60_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_60_BYTE_OFFSET = 13'h14a8;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_60_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_60_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_60_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_61_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_61_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_61_BYTE_OFFSET = 13'h14ac;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_61_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_61_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_61_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_62_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_62_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_62_BYTE_OFFSET = 13'h14b0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_62_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_62_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_62_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_63_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_63_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_63_BYTE_OFFSET = 13'h14b4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_63_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_63_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_63_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_64_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_64_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_64_BYTE_OFFSET = 13'h14b8;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_64_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_64_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_64_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_65_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_65_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_65_BYTE_OFFSET = 13'h14bc;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_65_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_65_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_65_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_66_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_66_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_66_BYTE_OFFSET = 13'h14c0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_66_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_66_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_66_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_67_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_67_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_67_BYTE_OFFSET = 13'h14c4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_67_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_67_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_67_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_68_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_68_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_68_BYTE_OFFSET = 13'h14c8;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_68_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_68_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_68_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_69_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_69_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_69_BYTE_OFFSET = 13'h14cc;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_69_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_69_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_69_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_70_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_70_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_70_BYTE_OFFSET = 13'h14d0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_70_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_70_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_70_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_71_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_71_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_71_BYTE_OFFSET = 13'h14d4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_71_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_71_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_71_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_72_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_72_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_72_BYTE_OFFSET = 13'h14d8;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_72_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_72_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_72_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_73_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_73_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_73_BYTE_OFFSET = 13'h14dc;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_73_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_73_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_73_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_74_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_74_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_74_BYTE_OFFSET = 13'h14e0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_74_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_74_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_74_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_75_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_75_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_75_BYTE_OFFSET = 13'h14e4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_75_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_75_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_75_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_76_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_76_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_76_BYTE_OFFSET = 13'h14e8;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_76_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_76_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_76_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_77_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_77_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_77_BYTE_OFFSET = 13'h14ec;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_77_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_77_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_77_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_78_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_78_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_78_BYTE_OFFSET = 13'h14f0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_78_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_78_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_78_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_79_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_79_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_79_BYTE_OFFSET = 13'h14f4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_79_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_79_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_79_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_80_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_80_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_80_BYTE_OFFSET = 13'h14f8;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_80_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_80_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_80_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_81_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_81_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_81_BYTE_OFFSET = 13'h14fc;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_81_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_81_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_81_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_82_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_82_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_82_BYTE_OFFSET = 13'h1500;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_82_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_82_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_82_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_83_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_83_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_83_BYTE_OFFSET = 13'h1504;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_83_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_83_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_83_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_84_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_84_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_84_BYTE_OFFSET = 13'h1508;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_84_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_84_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_84_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_85_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_85_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_85_BYTE_OFFSET = 13'h150c;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_85_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_85_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_85_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_86_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_86_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_86_BYTE_OFFSET = 13'h1510;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_86_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_86_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_86_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_87_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_87_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_87_BYTE_OFFSET = 13'h1514;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_87_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_87_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_87_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_88_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_88_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_88_BYTE_OFFSET = 13'h1518;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_88_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_88_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_88_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_89_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_89_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_89_BYTE_OFFSET = 13'h151c;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_89_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_89_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_89_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_90_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_90_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_90_BYTE_OFFSET = 13'h1520;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_90_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_90_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_90_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_91_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_91_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_91_BYTE_OFFSET = 13'h1524;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_91_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_91_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_91_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_92_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_92_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_92_BYTE_OFFSET = 13'h1528;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_92_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_92_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_92_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_93_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_93_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_93_BYTE_OFFSET = 13'h152c;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_93_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_93_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_93_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_94_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_94_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_94_BYTE_OFFSET = 13'h1530;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_94_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_94_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_94_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_95_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_95_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_95_BYTE_OFFSET = 13'h1534;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_95_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_95_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_95_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_96_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_96_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_96_BYTE_OFFSET = 13'h1538;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_96_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_96_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_96_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_97_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_97_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_97_BYTE_OFFSET = 13'h153c;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_97_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_97_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_97_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_98_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_98_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_98_BYTE_OFFSET = 13'h1540;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_98_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_98_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_98_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_99_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_99_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_99_BYTE_OFFSET = 13'h1544;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_99_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_99_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_99_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_100_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_100_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_100_BYTE_OFFSET = 13'h1548;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_100_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_100_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_100_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_101_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_101_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_101_BYTE_OFFSET = 13'h154c;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_101_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_101_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_101_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_102_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_102_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_102_BYTE_OFFSET = 13'h1550;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_102_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_102_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_102_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_103_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_103_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_103_BYTE_OFFSET = 13'h1554;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_103_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_103_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_103_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_104_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_104_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_104_BYTE_OFFSET = 13'h1558;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_104_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_104_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_104_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_105_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_105_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_105_BYTE_OFFSET = 13'h155c;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_105_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_105_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_105_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_106_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_106_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_106_BYTE_OFFSET = 13'h1560;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_106_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_106_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_106_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_107_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_107_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_107_BYTE_OFFSET = 13'h1564;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_107_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_107_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_107_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_108_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_108_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_108_BYTE_OFFSET = 13'h1568;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_108_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_108_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_108_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_109_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_109_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_109_BYTE_OFFSET = 13'h156c;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_109_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_109_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_109_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_110_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_110_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_110_BYTE_OFFSET = 13'h1570;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_110_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_110_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_110_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_111_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_111_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_111_BYTE_OFFSET = 13'h1574;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_111_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_111_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_111_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_112_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_112_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_112_BYTE_OFFSET = 13'h1578;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_112_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_112_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_112_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_113_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_113_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_113_BYTE_OFFSET = 13'h157c;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_113_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_113_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_113_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_114_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_114_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_114_BYTE_OFFSET = 13'h1580;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_114_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_114_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_114_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_115_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_115_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_115_BYTE_OFFSET = 13'h1584;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_115_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_115_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_115_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_116_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_116_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_116_BYTE_OFFSET = 13'h1588;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_116_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_116_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_116_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_117_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_117_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_117_BYTE_OFFSET = 13'h158c;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_117_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_117_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_117_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_118_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_118_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_118_BYTE_OFFSET = 13'h1590;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_118_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_118_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_118_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_119_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_119_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_119_BYTE_OFFSET = 13'h1594;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_119_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_119_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_119_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_120_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_120_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_120_BYTE_OFFSET = 13'h1598;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_120_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_120_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_120_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_121_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_121_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_121_BYTE_OFFSET = 13'h159c;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_121_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_121_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_121_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_122_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_122_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_122_BYTE_OFFSET = 13'h15a0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_122_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_122_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_122_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_123_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_123_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_123_BYTE_OFFSET = 13'h15a4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_123_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_123_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_123_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_124_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_124_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_124_BYTE_OFFSET = 13'h15a8;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_124_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_124_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_124_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_125_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_125_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_125_BYTE_OFFSET = 13'h15ac;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_125_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_125_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_125_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_126_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_126_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_126_BYTE_OFFSET = 13'h15b0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_126_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_126_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_126_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_127_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_127_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_127_BYTE_OFFSET = 13'h15b4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_127_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_127_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_127_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_128_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_128_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_128_BYTE_OFFSET = 13'h15b8;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_128_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_128_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_128_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_129_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_129_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_129_BYTE_OFFSET = 13'h15bc;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_129_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_129_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_129_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_130_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_130_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_130_BYTE_OFFSET = 13'h15c0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_130_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_130_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_130_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_131_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_131_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_131_BYTE_OFFSET = 13'h15c4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_131_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_131_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_131_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_132_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_132_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_132_BYTE_OFFSET = 13'h15c8;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_132_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_132_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_132_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_133_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_133_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_133_BYTE_OFFSET = 13'h15cc;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_133_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_133_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_133_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_134_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_134_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_134_BYTE_OFFSET = 13'h15d0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_134_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_134_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_134_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_135_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_135_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_135_BYTE_OFFSET = 13'h15d4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_135_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_135_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_135_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_136_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_136_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_136_BYTE_OFFSET = 13'h15d8;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_136_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_136_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_136_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_137_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_137_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_137_BYTE_OFFSET = 13'h15dc;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_137_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_137_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_137_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_138_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_138_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_138_BYTE_OFFSET = 13'h15e0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_138_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_138_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_138_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_139_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_139_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_139_BYTE_OFFSET = 13'h15e4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_139_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_139_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_139_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_140_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_140_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_140_BYTE_OFFSET = 13'h15e8;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_140_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_140_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_140_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_141_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_141_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_141_BYTE_OFFSET = 13'h15ec;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_141_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_141_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_141_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_142_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_142_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_142_BYTE_OFFSET = 13'h15f0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_142_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_142_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_142_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_143_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_143_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_143_BYTE_OFFSET = 13'h15f4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_143_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_143_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_143_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_144_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_144_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_144_BYTE_OFFSET = 13'h15f8;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_144_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_144_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_144_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_145_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_145_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_145_BYTE_OFFSET = 13'h15fc;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_145_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_145_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_145_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_146_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_146_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_146_BYTE_OFFSET = 13'h1600;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_146_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_146_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_146_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_147_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_147_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_147_BYTE_OFFSET = 13'h1604;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_147_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_147_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_147_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_148_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_148_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_148_BYTE_OFFSET = 13'h1608;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_148_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_148_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_148_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_149_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_149_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_149_BYTE_OFFSET = 13'h160c;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_149_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_149_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_149_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_150_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_150_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_150_BYTE_OFFSET = 13'h1610;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_150_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_150_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_150_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_151_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_151_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_151_BYTE_OFFSET = 13'h1614;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_151_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_151_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_151_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_152_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_152_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_152_BYTE_OFFSET = 13'h1618;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_152_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_152_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_152_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_153_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_153_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_153_BYTE_OFFSET = 13'h161c;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_153_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_153_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_153_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_154_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_154_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_154_BYTE_OFFSET = 13'h1620;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_154_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_154_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_154_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_155_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_155_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_155_BYTE_OFFSET = 13'h1624;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_155_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_155_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_155_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_156_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_156_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_156_BYTE_OFFSET = 13'h1628;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_156_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_156_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_156_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_157_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_157_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_157_BYTE_OFFSET = 13'h162c;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_157_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_157_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_157_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_158_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_158_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_158_BYTE_OFFSET = 13'h1630;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_158_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_158_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_158_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_159_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_159_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_159_BYTE_OFFSET = 13'h1634;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_159_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_159_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_159_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_160_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_160_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_160_BYTE_OFFSET = 13'h1638;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_160_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_160_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_160_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_161_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_161_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_161_BYTE_OFFSET = 13'h163c;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_161_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_161_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_161_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_162_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_162_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_162_BYTE_OFFSET = 13'h1640;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_162_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_162_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_162_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_163_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_163_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_163_BYTE_OFFSET = 13'h1644;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_163_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_163_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_163_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_164_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_164_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_164_BYTE_OFFSET = 13'h1648;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_164_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_164_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_164_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_165_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_165_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_165_BYTE_OFFSET = 13'h164c;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_165_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_165_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_165_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_166_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_166_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_166_BYTE_OFFSET = 13'h1650;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_166_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_166_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_166_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_167_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_167_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_167_BYTE_OFFSET = 13'h1654;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_167_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_167_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_167_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_168_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_168_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_168_BYTE_OFFSET = 13'h1658;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_168_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_168_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_168_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_169_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_169_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_169_BYTE_OFFSET = 13'h165c;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_169_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_169_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_169_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_170_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_170_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_170_BYTE_OFFSET = 13'h1660;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_170_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_170_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_170_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_171_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_171_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_171_BYTE_OFFSET = 13'h1664;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_171_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_171_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_171_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_172_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_172_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_172_BYTE_OFFSET = 13'h1668;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_172_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_172_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_172_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_173_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_173_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_173_BYTE_OFFSET = 13'h166c;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_173_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_173_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_173_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_174_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_174_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_174_BYTE_OFFSET = 13'h1670;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_174_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_174_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_174_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_175_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_175_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_175_BYTE_OFFSET = 13'h1674;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_175_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_175_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_175_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_176_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_176_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_176_BYTE_OFFSET = 13'h1678;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_176_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_176_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_176_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_177_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_177_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_177_BYTE_OFFSET = 13'h167c;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_177_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_177_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_177_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_178_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_178_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_178_BYTE_OFFSET = 13'h1680;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_178_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_178_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_178_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_179_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_179_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_179_BYTE_OFFSET = 13'h1684;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_179_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_179_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_179_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_180_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_180_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_180_BYTE_OFFSET = 13'h1688;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_180_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_180_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_180_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_181_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_181_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_181_BYTE_OFFSET = 13'h168c;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_181_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_181_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_181_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_182_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_182_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_182_BYTE_OFFSET = 13'h1690;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_182_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_182_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_182_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_183_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_183_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_183_BYTE_OFFSET = 13'h1694;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_183_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_183_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_183_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_184_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_184_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_184_BYTE_OFFSET = 13'h1698;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_184_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_184_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_184_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_185_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_185_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_185_BYTE_OFFSET = 13'h169c;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_185_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_185_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_185_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_186_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_186_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_186_BYTE_OFFSET = 13'h16a0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_186_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_186_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_186_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_187_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_187_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_187_BYTE_OFFSET = 13'h16a4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_187_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_187_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_187_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_188_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_188_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_188_BYTE_OFFSET = 13'h16a8;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_188_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_188_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_188_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_189_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_189_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_189_BYTE_OFFSET = 13'h16ac;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_189_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_189_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_189_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_190_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_190_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_190_BYTE_OFFSET = 13'h16b0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_190_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_190_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_190_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_191_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_191_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_191_BYTE_OFFSET = 13'h16b4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_191_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_191_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_191_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_192_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_192_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_192_BYTE_OFFSET = 13'h16b8;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_192_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_192_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_192_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_193_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_193_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_193_BYTE_OFFSET = 13'h16bc;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_193_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_193_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_193_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_194_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_194_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_194_BYTE_OFFSET = 13'h16c0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_194_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_194_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_194_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_195_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_195_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_195_BYTE_OFFSET = 13'h16c4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_195_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_195_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_195_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_196_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_196_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_196_BYTE_OFFSET = 13'h16c8;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_196_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_196_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_196_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_197_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_197_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_197_BYTE_OFFSET = 13'h16cc;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_197_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_197_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_197_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_198_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_198_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_198_BYTE_OFFSET = 13'h16d0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_198_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_198_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_198_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_199_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_199_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_199_BYTE_OFFSET = 13'h16d4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_199_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_199_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_199_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_200_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_200_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_200_BYTE_OFFSET = 13'h16d8;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_200_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_200_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_200_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_201_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_201_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_201_BYTE_OFFSET = 13'h16dc;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_201_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_201_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_201_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_202_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_202_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_202_BYTE_OFFSET = 13'h16e0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_202_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_202_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_202_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_203_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_203_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_203_BYTE_OFFSET = 13'h16e4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_203_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_203_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_203_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_204_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_204_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_204_BYTE_OFFSET = 13'h16e8;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_204_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_204_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_204_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_205_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_205_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_205_BYTE_OFFSET = 13'h16ec;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_205_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_205_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_205_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_206_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_206_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_206_BYTE_OFFSET = 13'h16f0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_206_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_206_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_206_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_207_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_207_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_CODEWRD_OUT_BIT_207_BYTE_OFFSET = 13'h16f4;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_207_FINAL_CWORD_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_CODEWRD_OUT_BIT_207_FINAL_CWORD_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_CODEWRD_OUT_BIT_207_FINAL_CWORD_BIT_OFFSET = 0;
  localparam int LDPC_DEC_PASS_FAIL_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_PASS_FAIL_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_PASS_FAIL_BYTE_OFFSET = 13'h16f8;
  localparam int LDPC_DEC_PASS_FAIL_PASS_FAIL_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_PASS_FAIL_PASS_FAIL_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_PASS_FAIL_PASS_FAIL_BIT_OFFSET = 0;
  localparam int LDPC_DEC_PASS_FAIL_DECODER_BYTE_WIDTH = 4;
  localparam int LDPC_DEC_PASS_FAIL_DECODER_BYTE_SIZE = 4;
  localparam bit [12:0] LDPC_DEC_PASS_FAIL_DECODER_BYTE_OFFSET = 13'h16fc;
  localparam int LDPC_DEC_PASS_FAIL_DECODER_PASS_FAIL_DECODER_BIT_BIT_WIDTH = 1;
  localparam bit LDPC_DEC_PASS_FAIL_DECODER_PASS_FAIL_DECODER_BIT_BIT_MASK = 1'h1;
  localparam int LDPC_DEC_PASS_FAIL_DECODER_PASS_FAIL_DECODER_BIT_BIT_OFFSET = 0;
endpackage
