              flogtanh0x00002_0 = 
          (!flogtanh_sel[1]) ? 
                       flogtanh0x00001_0_q: 
                       flogtanh0x00001_1_q;
              flogtanh0x00002_1 = 
          (!flogtanh_sel[1]) ? 
                       flogtanh0x00001_2_q: 
                       flogtanh0x00001_3_q;
              flogtanh0x00002_2 = 
          (!flogtanh_sel[1]) ? 
                       flogtanh0x00001_4_q: 
                       flogtanh0x00001_5_q;
              flogtanh0x00002_3 = 
          (!flogtanh_sel[1]) ? 
                       flogtanh0x00001_6_q: 
                       flogtanh0x00001_7_q;
              flogtanh0x00002_4 = 
          (!flogtanh_sel[1]) ? 
                       flogtanh0x00001_8_q: 
                       flogtanh0x00001_9_q;
              flogtanh0x00002_5 = 
          (!flogtanh_sel[1]) ? 
                       flogtanh0x00001_10_q: 
                       flogtanh0x00001_11_q;
              flogtanh0x00002_6 = 
          (!flogtanh_sel[1]) ? 
                       flogtanh0x00001_12_q: 
                       flogtanh0x00001_13_q;
              flogtanh0x00002_7 = 
          (!flogtanh_sel[1]) ? 
                       flogtanh0x00001_14_q: 
                       flogtanh0x00001_15_q;
              flogtanh0x00002_8 = 
          (!flogtanh_sel[1]) ? 
                       flogtanh0x00001_16_q: 
                       flogtanh0x00001_17_q;
              flogtanh0x00002_9 = 
          (!flogtanh_sel[1]) ? 
                       flogtanh0x00001_18_q: 
                       flogtanh0x00001_19_q;
              flogtanh0x00002_10 = 
          (!flogtanh_sel[1]) ? 
                       flogtanh0x00001_20_q: 
                       flogtanh0x00001_21_q;
              flogtanh0x00002_11 = 
          (!flogtanh_sel[1]) ? 
                       flogtanh0x00001_22_q: 
                       flogtanh0x00001_23_q;
              flogtanh0x00002_12 = 
          (!flogtanh_sel[1]) ? 
                       flogtanh0x00001_24_q: 
                       flogtanh0x00001_25_q;
              flogtanh0x00002_13 = 
          (!flogtanh_sel[1]) ? 
                       flogtanh0x00001_26_q: 
                       flogtanh0x00001_27_q;
              flogtanh0x00002_14 = 
          (!flogtanh_sel[1]) ? 
                       flogtanh0x00001_28_q: 
                       flogtanh0x00001_29_q;
              flogtanh0x00002_15 = 
          (!flogtanh_sel[1]) ? 
                       flogtanh0x00001_30_q: 
                       flogtanh0x00001_31_q;
              flogtanh0x00002_16 = 
          (!flogtanh_sel[1]) ? 
                       flogtanh0x00001_32_q: 
                       flogtanh0x00001_33_q;
              flogtanh0x00002_17 = 
          (!flogtanh_sel[1]) ? 
                       flogtanh0x00001_34_q: 
                       flogtanh0x00001_35_q;
              flogtanh0x00002_18 = 
          (!flogtanh_sel[1]) ? 
                       flogtanh0x00001_36_q: 
                       flogtanh0x00001_37_q;
              flogtanh0x00002_19 = 
          (!flogtanh_sel[1]) ? 
                       flogtanh0x00001_38_q: 
                       flogtanh0x00001_39_q;
              flogtanh0x00002_20 = 
          (!flogtanh_sel[1]) ? 
                       flogtanh0x00001_40_q: 
                       flogtanh0x00001_41_q;
              flogtanh0x00002_21 = 
          (!flogtanh_sel[1]) ? 
                       flogtanh0x00001_42_q: 
                       flogtanh0x00001_43_q;
              flogtanh0x00002_22 = 
          (!flogtanh_sel[1]) ? 
                       flogtanh0x00001_44_q: 
                       flogtanh0x00001_45_q;
              flogtanh0x00002_23 = 
          (!flogtanh_sel[1]) ? 
                       flogtanh0x00001_46_q: 
                       flogtanh0x00001_47_q;
              flogtanh0x00002_24 = 
          (!flogtanh_sel[1]) ? 
                       flogtanh0x00001_48_q: 
                       flogtanh0x00001_49_q;
              flogtanh0x00002_25 = 
          (!flogtanh_sel[1]) ? 
                       flogtanh0x00001_50_q: 
                       flogtanh0x00001_51_q;
              flogtanh0x00002_26 = 
          (!flogtanh_sel[1]) ? 
                       flogtanh0x00001_52_q: 
                       flogtanh0x00001_53_q;
              flogtanh0x00002_27 = 
          (!flogtanh_sel[1]) ? 
                       flogtanh0x00001_54_q: 
                       flogtanh0x00001_55_q;
              flogtanh0x00002_28 = 
          (!flogtanh_sel[1]) ? 
                       flogtanh0x00001_56_q: 
                       flogtanh0x00001_57_q;
              flogtanh0x00002_29 = 
          (!flogtanh_sel[1]) ? 
                       flogtanh0x00001_58_q: 
                       flogtanh0x00001_59_q;
              flogtanh0x00002_30 = 
          (!flogtanh_sel[1]) ? 
                       flogtanh0x00001_60_q: 
                       flogtanh0x00001_61_q;
              flogtanh0x00002_31 = 
          (!flogtanh_sel[1]) ? 
                       flogtanh0x00001_62_q: 
                       flogtanh0x00001_63_q;
               flogtanh0x00002_32 =  flogtanh0x00001_64_q ;
               flogtanh0x00002_33 =  flogtanh0x00001_66_q ;
               flogtanh0x00002_34 =  flogtanh0x00001_68_q ;
               flogtanh0x00002_35 =  flogtanh0x00001_70_q ;
              flogtanh0x00002_36 = 
          (!flogtanh_sel[1]) ? 
                       flogtanh0x00001_72_q: 
                       flogtanh0x00001_73_q;
              flogtanh0x00002_37 = 
          (!flogtanh_sel[1]) ? 
                       flogtanh0x00001_74_q: 
                       flogtanh0x00001_75_q;
              flogtanh0x00002_38 = 
          (!flogtanh_sel[1]) ? 
                       flogtanh0x00001_76_q: 
                       flogtanh0x00001_77_q;
               flogtanh0x00002_39 =  flogtanh0x00001_78_q ;
              flogtanh0x00002_40 = 
          (!flogtanh_sel[1]) ? 
                       flogtanh0x00001_80_q: 
                       flogtanh0x00001_81_q;
              flogtanh0x00002_41 = 
          (!flogtanh_sel[1]) ? 
                       flogtanh0x00001_82_q: 
                       flogtanh0x00001_83_q;
               flogtanh0x00002_42 =  flogtanh0x00001_84_q ;
              flogtanh0x00002_43 = 
          (!flogtanh_sel[1]) ? 
                       flogtanh0x00001_86_q: 
                       flogtanh0x00001_87_q;
               flogtanh0x00002_44 =  flogtanh0x00001_88_q ;
              flogtanh0x00002_45 = 
          (!flogtanh_sel[1]) ? 
                       flogtanh0x00001_90_q: 
                       flogtanh0x00001_91_q;
               flogtanh0x00002_46 =  flogtanh0x00001_92_q ;
              flogtanh0x00002_47 = 
          (!flogtanh_sel[1]) ? 
                       flogtanh0x00001_94_q: 
                       flogtanh0x00001_95_q;
               flogtanh0x00002_48 =  flogtanh0x00001_96_q ;
               flogtanh0x00002_49 =  flogtanh0x00001_98_q ;
              flogtanh0x00002_50 = 
          (!flogtanh_sel[1]) ? 
                       flogtanh0x00001_100_q: 
                       flogtanh0x00001_101_q;
               flogtanh0x00002_51 =  flogtanh0x00001_102_q ;
               flogtanh0x00002_52 =  flogtanh0x00001_104_q ;
              flogtanh0x00002_53 = 
          (!flogtanh_sel[1]) ? 
                       flogtanh0x00001_106_q: 
                       flogtanh0x00001_107_q;
               flogtanh0x00002_54 =  flogtanh0x00001_108_q ;
               flogtanh0x00002_55 =  flogtanh0x00001_110_q ;
               flogtanh0x00002_56 =  flogtanh0x00001_112_q ;
              flogtanh0x00002_57 = 
          (!flogtanh_sel[1]) ? 
                       flogtanh0x00001_114_q: 
                       flogtanh0x00001_115_q;
               flogtanh0x00002_58 =  flogtanh0x00001_116_q ;
               flogtanh0x00002_59 =  flogtanh0x00001_118_q ;
               flogtanh0x00002_60 =  flogtanh0x00001_120_q ;
               flogtanh0x00002_61 =  flogtanh0x00001_122_q ;
               flogtanh0x00002_62 =  flogtanh0x00001_124_q ;
               flogtanh0x00002_63 =  flogtanh0x00001_126_q ;
               flogtanh0x00002_64 =  flogtanh0x00001_128_q ;
               flogtanh0x00002_65 =  flogtanh0x00001_130_q ;
               flogtanh0x00002_66 =  flogtanh0x00001_132_q ;
               flogtanh0x00002_67 =  flogtanh0x00001_134_q ;
               flogtanh0x00002_68 =  flogtanh0x00001_136_q ;
               flogtanh0x00002_69 =  flogtanh0x00001_138_q ;
               flogtanh0x00002_70 =  flogtanh0x00001_140_q ;
              flogtanh0x00002_71 = 
          (!flogtanh_sel[1]) ? 
                       flogtanh0x00001_142_q: 
                       flogtanh0x00001_143_q;
               flogtanh0x00002_72 =  flogtanh0x00001_144_q ;
               flogtanh0x00002_73 =  flogtanh0x00001_146_q ;
               flogtanh0x00002_74 =  flogtanh0x00001_148_q ;
               flogtanh0x00002_75 =  flogtanh0x00001_150_q ;
               flogtanh0x00002_76 =  flogtanh0x00001_152_q ;
               flogtanh0x00002_77 =  flogtanh0x00001_154_q ;
               flogtanh0x00002_78 =  flogtanh0x00001_156_q ;
               flogtanh0x00002_79 =  flogtanh0x00001_158_q ;
               flogtanh0x00002_80 =  flogtanh0x00001_160_q ;
               flogtanh0x00002_81 =  flogtanh0x00001_162_q ;
               flogtanh0x00002_82 =  flogtanh0x00001_164_q ;
               flogtanh0x00002_83 =  flogtanh0x00001_166_q ;
               flogtanh0x00002_84 =  flogtanh0x00001_168_q ;
               flogtanh0x00002_85 =  flogtanh0x00001_170_q ;
               flogtanh0x00002_86 =  flogtanh0x00001_172_q ;
               flogtanh0x00002_87 =  flogtanh0x00001_174_q ;
              flogtanh0x00002_88 = 
          (!flogtanh_sel[1]) ? 
                       flogtanh0x00001_176_q: 
                       flogtanh0x00001_177_q;
               flogtanh0x00002_89 =  0;
