reg [flogtanh_WDTH -1:0] flogtanh0x00004_0, flogtanh0x00004_0_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00004_1, flogtanh0x00004_1_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00004_2, flogtanh0x00004_2_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00004_3, flogtanh0x00004_3_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00004_4, flogtanh0x00004_4_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00004_5, flogtanh0x00004_5_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00004_6, flogtanh0x00004_6_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00004_7, flogtanh0x00004_7_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00004_8, flogtanh0x00004_8_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00004_9, flogtanh0x00004_9_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00004_10, flogtanh0x00004_10_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00004_11, flogtanh0x00004_11_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00004_12, flogtanh0x00004_12_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00004_13, flogtanh0x00004_13_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00004_14, flogtanh0x00004_14_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00004_15, flogtanh0x00004_15_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00004_16, flogtanh0x00004_16_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00004_17, flogtanh0x00004_17_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00004_18, flogtanh0x00004_18_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00004_19, flogtanh0x00004_19_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00004_20, flogtanh0x00004_20_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00004_21, flogtanh0x00004_21_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00004_22, flogtanh0x00004_22_q;
reg [flogtanh_WDTH -1:0] flogtanh0x00004_23, flogtanh0x00004_23_q;
reg start_d_flogtanh0x00004_q ;
always_comb begin
 flogtanh0x00004_0_q =  flogtanh0x00004_0;
 flogtanh0x00004_1_q =  flogtanh0x00004_1;
 flogtanh0x00004_2_q =  flogtanh0x00004_2;
 flogtanh0x00004_3_q =  flogtanh0x00004_3;
 flogtanh0x00004_4_q =  flogtanh0x00004_4;
 flogtanh0x00004_5_q =  flogtanh0x00004_5;
 flogtanh0x00004_6_q =  flogtanh0x00004_6;
 flogtanh0x00004_7_q =  flogtanh0x00004_7;
 flogtanh0x00004_8_q =  flogtanh0x00004_8;
 flogtanh0x00004_9_q =  flogtanh0x00004_9;
 flogtanh0x00004_10_q =  flogtanh0x00004_10;
 flogtanh0x00004_11_q =  flogtanh0x00004_11;
 flogtanh0x00004_12_q =  flogtanh0x00004_12;
 flogtanh0x00004_13_q =  flogtanh0x00004_13;
 flogtanh0x00004_14_q =  flogtanh0x00004_14;
 flogtanh0x00004_15_q =  flogtanh0x00004_15;
 flogtanh0x00004_16_q =  flogtanh0x00004_16;
 flogtanh0x00004_17_q =  flogtanh0x00004_17;
 flogtanh0x00004_18_q =  flogtanh0x00004_18;
 flogtanh0x00004_19_q =  flogtanh0x00004_19;
 flogtanh0x00004_20_q =  flogtanh0x00004_20;
 flogtanh0x00004_21_q =  flogtanh0x00004_21;
 flogtanh0x00004_22_q =  flogtanh0x00004_22;
 flogtanh0x00004_23_q =  flogtanh0x00004_23;
 start_d_flogtanh0x00004_q =  start_d_flogtanh0x00003_q;
end
