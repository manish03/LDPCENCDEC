`define SIM_RAM 1
