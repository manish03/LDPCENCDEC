              flogtanh0x00006_0 = 
          (!flogtanh_sel[5]) ? 
                       flogtanh0x00005_0_q: 
                       flogtanh0x00005_1_q;
              flogtanh0x00006_1 = 
          (!flogtanh_sel[5]) ? 
                       flogtanh0x00005_2_q: 
                       flogtanh0x00005_3_q;
              flogtanh0x00006_2 = 
          (!flogtanh_sel[5]) ? 
                       flogtanh0x00005_4_q: 
                       flogtanh0x00005_5_q;
              flogtanh0x00006_3 = 
          (!flogtanh_sel[5]) ? 
                       flogtanh0x00005_6_q: 
                       flogtanh0x00005_7_q;
              flogtanh0x00006_4 = 
          (!flogtanh_sel[5]) ? 
                       flogtanh0x00005_8_q: 
                       flogtanh0x00005_9_q;
              flogtanh0x00006_5 = 
          (!flogtanh_sel[5]) ? 
                       flogtanh0x00005_10_q: 
                       flogtanh0x00005_11_q;
