              flogtanh0x00004_0 = 
          (!flogtanh_sel[3]) ? 
                       flogtanh0x00003_0_q: 
                       flogtanh0x00003_1_q;
              flogtanh0x00004_1 = 
          (!flogtanh_sel[3]) ? 
                       flogtanh0x00003_2_q: 
                       flogtanh0x00003_3_q;
              flogtanh0x00004_2 = 
          (!flogtanh_sel[3]) ? 
                       flogtanh0x00003_4_q: 
                       flogtanh0x00003_5_q;
              flogtanh0x00004_3 = 
          (!flogtanh_sel[3]) ? 
                       flogtanh0x00003_6_q: 
                       flogtanh0x00003_7_q;
              flogtanh0x00004_4 = 
          (!flogtanh_sel[3]) ? 
                       flogtanh0x00003_8_q: 
                       flogtanh0x00003_9_q;
              flogtanh0x00004_5 = 
          (!flogtanh_sel[3]) ? 
                       flogtanh0x00003_10_q: 
                       flogtanh0x00003_11_q;
              flogtanh0x00004_6 = 
          (!flogtanh_sel[3]) ? 
                       flogtanh0x00003_12_q: 
                       flogtanh0x00003_13_q;
              flogtanh0x00004_7 = 
          (!flogtanh_sel[3]) ? 
                       flogtanh0x00003_14_q: 
                       flogtanh0x00003_15_q;
              flogtanh0x00004_8 = 
          (!flogtanh_sel[3]) ? 
                       flogtanh0x00003_16_q: 
                       flogtanh0x00003_17_q;
              flogtanh0x00004_9 = 
          (!flogtanh_sel[3]) ? 
                       flogtanh0x00003_18_q: 
                       flogtanh0x00003_19_q;
              flogtanh0x00004_10 = 
          (!flogtanh_sel[3]) ? 
                       flogtanh0x00003_20_q: 
                       flogtanh0x00003_21_q;
              flogtanh0x00004_11 = 
          (!flogtanh_sel[3]) ? 
                       flogtanh0x00003_22_q: 
                       flogtanh0x00003_23_q;
              flogtanh0x00004_12 = 
          (!flogtanh_sel[3]) ? 
                       flogtanh0x00003_24_q: 
                       flogtanh0x00003_25_q;
              flogtanh0x00004_13 = 
          (!flogtanh_sel[3]) ? 
                       flogtanh0x00003_26_q: 
                       flogtanh0x00003_27_q;
              flogtanh0x00004_14 = 
          (!flogtanh_sel[3]) ? 
                       flogtanh0x00003_28_q: 
                       flogtanh0x00003_29_q;
              flogtanh0x00004_15 = 
          (!flogtanh_sel[3]) ? 
                       flogtanh0x00003_30_q: 
                       flogtanh0x00003_31_q;
               flogtanh0x00004_16 =  flogtanh0x00003_32_q ;
              flogtanh0x00004_17 = 
          (!flogtanh_sel[3]) ? 
                       flogtanh0x00003_34_q: 
                       flogtanh0x00003_35_q;
               flogtanh0x00004_18 =  flogtanh0x00003_36_q ;
               flogtanh0x00004_19 =  flogtanh0x00003_38_q ;
               flogtanh0x00004_20 =  flogtanh0x00003_40_q ;
               flogtanh0x00004_21 =  flogtanh0x00003_42_q ;
              flogtanh0x00004_22 = 
          (!flogtanh_sel[3]) ? 
                       flogtanh0x00003_44_q: 
                       flogtanh0x00003_45_q;
               flogtanh0x00004_23 =  0;
