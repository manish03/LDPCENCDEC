wire o_LDPC_ENC_MSG_IN_0_msg_in;
wire o_LDPC_ENC_MSG_IN_1_msg_in;
wire o_LDPC_ENC_MSG_IN_2_msg_in;
wire o_LDPC_ENC_MSG_IN_3_msg_in;
wire o_LDPC_ENC_MSG_IN_4_msg_in;
wire o_LDPC_ENC_MSG_IN_5_msg_in;
wire o_LDPC_ENC_MSG_IN_6_msg_in;
wire o_LDPC_ENC_MSG_IN_7_msg_in;
wire o_LDPC_ENC_MSG_IN_8_msg_in;
wire o_LDPC_ENC_MSG_IN_9_msg_in;
wire o_LDPC_ENC_MSG_IN_10_msg_in;
wire o_LDPC_ENC_MSG_IN_11_msg_in;
wire o_LDPC_ENC_MSG_IN_12_msg_in;
wire o_LDPC_ENC_MSG_IN_13_msg_in;
wire o_LDPC_ENC_MSG_IN_14_msg_in;
wire o_LDPC_ENC_MSG_IN_15_msg_in;
wire o_LDPC_ENC_MSG_IN_16_msg_in;
wire o_LDPC_ENC_MSG_IN_17_msg_in;
wire o_LDPC_ENC_MSG_IN_18_msg_in;
wire o_LDPC_ENC_MSG_IN_19_msg_in;
wire o_LDPC_ENC_MSG_IN_20_msg_in;
wire o_LDPC_ENC_MSG_IN_21_msg_in;
wire o_LDPC_ENC_MSG_IN_22_msg_in;
wire o_LDPC_ENC_MSG_IN_23_msg_in;
wire o_LDPC_ENC_MSG_IN_24_msg_in;
wire o_LDPC_ENC_MSG_IN_25_msg_in;
wire o_LDPC_ENC_MSG_IN_26_msg_in;
wire o_LDPC_ENC_MSG_IN_27_msg_in;
wire o_LDPC_ENC_MSG_IN_28_msg_in;
wire o_LDPC_ENC_MSG_IN_29_msg_in;
wire o_LDPC_ENC_MSG_IN_30_msg_in;
wire o_LDPC_ENC_MSG_IN_31_msg_in;
wire o_LDPC_ENC_MSG_IN_32_msg_in;
wire o_LDPC_ENC_MSG_IN_33_msg_in;
wire o_LDPC_ENC_MSG_IN_34_msg_in;
wire o_LDPC_ENC_MSG_IN_35_msg_in;
wire o_LDPC_ENC_MSG_IN_36_msg_in;
wire o_LDPC_ENC_MSG_IN_37_msg_in;
wire o_LDPC_ENC_MSG_IN_38_msg_in;
wire o_LDPC_ENC_MSG_IN_39_msg_in;
wire i_LDPC_ENC_CODEWRD_OUT_0_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_1_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_2_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_3_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_4_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_5_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_6_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_7_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_8_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_9_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_10_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_11_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_12_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_13_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_14_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_15_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_16_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_17_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_18_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_19_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_20_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_21_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_22_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_23_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_24_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_25_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_26_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_27_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_28_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_29_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_30_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_31_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_32_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_33_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_34_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_35_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_36_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_37_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_38_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_39_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_40_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_41_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_42_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_43_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_44_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_45_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_46_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_47_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_48_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_49_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_50_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_51_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_52_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_53_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_54_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_55_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_56_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_57_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_58_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_59_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_60_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_61_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_62_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_63_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_64_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_65_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_66_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_67_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_68_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_69_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_70_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_71_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_72_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_73_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_74_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_75_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_76_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_77_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_78_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_79_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_80_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_81_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_82_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_83_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_84_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_85_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_86_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_87_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_88_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_89_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_90_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_91_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_92_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_93_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_94_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_95_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_96_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_97_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_98_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_99_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_100_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_101_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_102_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_103_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_104_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_105_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_106_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_107_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_108_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_109_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_110_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_111_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_112_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_113_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_114_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_115_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_116_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_117_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_118_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_119_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_120_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_121_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_122_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_123_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_124_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_125_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_126_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_127_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_128_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_129_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_130_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_131_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_132_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_133_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_134_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_135_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_136_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_137_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_138_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_139_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_140_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_141_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_142_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_143_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_144_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_145_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_146_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_147_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_148_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_149_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_150_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_151_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_152_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_153_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_154_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_155_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_156_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_157_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_158_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_159_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_160_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_161_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_162_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_163_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_164_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_165_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_166_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_167_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_168_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_169_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_170_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_171_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_172_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_173_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_174_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_175_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_176_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_177_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_178_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_179_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_180_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_181_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_182_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_183_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_184_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_185_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_186_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_187_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_188_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_189_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_190_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_191_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_192_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_193_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_194_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_195_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_196_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_197_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_198_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_199_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_200_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_201_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_202_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_203_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_204_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_205_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_206_enc_codeword;
wire i_LDPC_ENC_CODEWRD_OUT_207_enc_codeword;
wire i_LDPC_ENC_CODEWRD_VLD_enc_codeword_valid;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_0_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_1_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_2_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_3_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_4_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_5_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_6_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_7_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_8_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_9_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_10_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_11_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_12_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_13_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_14_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_15_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_16_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_17_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_18_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_19_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_20_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_21_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_22_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_23_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_24_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_25_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_26_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_27_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_28_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_29_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_30_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_31_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_32_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_33_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_34_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_35_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_36_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_37_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_38_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_39_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_40_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_41_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_42_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_43_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_44_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_45_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_46_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_47_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_48_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_49_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_50_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_51_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_52_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_53_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_54_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_55_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_56_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_57_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_58_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_59_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_60_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_61_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_62_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_63_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_64_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_65_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_66_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_67_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_68_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_69_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_70_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_71_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_72_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_73_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_74_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_75_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_76_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_77_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_78_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_79_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_80_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_81_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_82_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_83_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_84_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_85_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_86_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_87_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_88_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_89_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_90_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_91_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_92_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_93_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_94_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_95_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_96_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_97_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_98_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_99_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_100_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_101_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_102_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_103_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_104_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_105_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_106_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_107_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_108_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_109_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_110_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_111_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_112_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_113_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_114_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_115_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_116_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_117_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_118_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_119_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_120_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_121_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_122_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_123_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_124_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_125_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_126_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_127_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_128_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_129_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_130_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_131_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_132_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_133_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_134_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_135_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_136_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_137_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_138_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_139_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_140_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_141_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_142_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_143_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_144_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_145_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_146_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_147_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_148_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_149_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_150_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_151_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_152_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_153_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_154_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_155_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_156_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_157_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_158_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_159_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_160_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_161_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_162_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_163_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_164_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_165_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_166_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_167_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_168_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_169_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_170_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_171_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_172_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_173_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_174_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_175_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_176_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_177_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_178_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_179_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_180_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_181_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_182_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_183_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_184_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_185_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_186_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_187_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_188_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_189_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_190_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_191_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_192_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_193_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_194_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_195_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_196_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_197_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_198_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_199_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_200_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_201_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_202_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_203_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_204_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_205_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_206_cword_q0;
wire [1:0] o_LDPC_DEC_CODEWRD_IN_207_cword_q0;
wire o_LDPC_DEC_ERR_INTRODUCED_err_intro;
wire o_LDPC_DEC_EXPSYND_0_exp_syn;
wire o_LDPC_DEC_EXPSYND_1_exp_syn;
wire o_LDPC_DEC_EXPSYND_2_exp_syn;
wire o_LDPC_DEC_EXPSYND_3_exp_syn;
wire o_LDPC_DEC_EXPSYND_4_exp_syn;
wire o_LDPC_DEC_EXPSYND_5_exp_syn;
wire o_LDPC_DEC_EXPSYND_6_exp_syn;
wire o_LDPC_DEC_EXPSYND_7_exp_syn;
wire o_LDPC_DEC_EXPSYND_8_exp_syn;
wire o_LDPC_DEC_EXPSYND_9_exp_syn;
wire o_LDPC_DEC_EXPSYND_10_exp_syn;
wire o_LDPC_DEC_EXPSYND_11_exp_syn;
wire o_LDPC_DEC_EXPSYND_12_exp_syn;
wire o_LDPC_DEC_EXPSYND_13_exp_syn;
wire o_LDPC_DEC_EXPSYND_14_exp_syn;
wire o_LDPC_DEC_EXPSYND_15_exp_syn;
wire o_LDPC_DEC_EXPSYND_16_exp_syn;
wire o_LDPC_DEC_EXPSYND_17_exp_syn;
wire o_LDPC_DEC_EXPSYND_18_exp_syn;
wire o_LDPC_DEC_EXPSYND_19_exp_syn;
wire o_LDPC_DEC_EXPSYND_20_exp_syn;
wire o_LDPC_DEC_EXPSYND_21_exp_syn;
wire o_LDPC_DEC_EXPSYND_22_exp_syn;
wire o_LDPC_DEC_EXPSYND_23_exp_syn;
wire o_LDPC_DEC_EXPSYND_24_exp_syn;
wire o_LDPC_DEC_EXPSYND_25_exp_syn;
wire o_LDPC_DEC_EXPSYND_26_exp_syn;
wire o_LDPC_DEC_EXPSYND_27_exp_syn;
wire o_LDPC_DEC_EXPSYND_28_exp_syn;
wire o_LDPC_DEC_EXPSYND_29_exp_syn;
wire o_LDPC_DEC_EXPSYND_30_exp_syn;
wire o_LDPC_DEC_EXPSYND_31_exp_syn;
wire o_LDPC_DEC_EXPSYND_32_exp_syn;
wire o_LDPC_DEC_EXPSYND_33_exp_syn;
wire o_LDPC_DEC_EXPSYND_34_exp_syn;
wire o_LDPC_DEC_EXPSYND_35_exp_syn;
wire o_LDPC_DEC_EXPSYND_36_exp_syn;
wire o_LDPC_DEC_EXPSYND_37_exp_syn;
wire o_LDPC_DEC_EXPSYND_38_exp_syn;
wire o_LDPC_DEC_EXPSYND_39_exp_syn;
wire o_LDPC_DEC_EXPSYND_40_exp_syn;
wire o_LDPC_DEC_EXPSYND_41_exp_syn;
wire o_LDPC_DEC_EXPSYND_42_exp_syn;
wire o_LDPC_DEC_EXPSYND_43_exp_syn;
wire o_LDPC_DEC_EXPSYND_44_exp_syn;
wire o_LDPC_DEC_EXPSYND_45_exp_syn;
wire o_LDPC_DEC_EXPSYND_46_exp_syn;
wire o_LDPC_DEC_EXPSYND_47_exp_syn;
wire o_LDPC_DEC_EXPSYND_48_exp_syn;
wire o_LDPC_DEC_EXPSYND_49_exp_syn;
wire o_LDPC_DEC_EXPSYND_50_exp_syn;
wire o_LDPC_DEC_EXPSYND_51_exp_syn;
wire o_LDPC_DEC_EXPSYND_52_exp_syn;
wire o_LDPC_DEC_EXPSYND_53_exp_syn;
wire o_LDPC_DEC_EXPSYND_54_exp_syn;
wire o_LDPC_DEC_EXPSYND_55_exp_syn;
wire o_LDPC_DEC_EXPSYND_56_exp_syn;
wire o_LDPC_DEC_EXPSYND_57_exp_syn;
wire o_LDPC_DEC_EXPSYND_58_exp_syn;
wire o_LDPC_DEC_EXPSYND_59_exp_syn;
wire o_LDPC_DEC_EXPSYND_60_exp_syn;
wire o_LDPC_DEC_EXPSYND_61_exp_syn;
wire o_LDPC_DEC_EXPSYND_62_exp_syn;
wire o_LDPC_DEC_EXPSYND_63_exp_syn;
wire o_LDPC_DEC_EXPSYND_64_exp_syn;
wire o_LDPC_DEC_EXPSYND_65_exp_syn;
wire o_LDPC_DEC_EXPSYND_66_exp_syn;
wire o_LDPC_DEC_EXPSYND_67_exp_syn;
wire o_LDPC_DEC_EXPSYND_68_exp_syn;
wire o_LDPC_DEC_EXPSYND_69_exp_syn;
wire o_LDPC_DEC_EXPSYND_70_exp_syn;
wire o_LDPC_DEC_EXPSYND_71_exp_syn;
wire o_LDPC_DEC_EXPSYND_72_exp_syn;
wire o_LDPC_DEC_EXPSYND_73_exp_syn;
wire o_LDPC_DEC_EXPSYND_74_exp_syn;
wire o_LDPC_DEC_EXPSYND_75_exp_syn;
wire o_LDPC_DEC_EXPSYND_76_exp_syn;
wire o_LDPC_DEC_EXPSYND_77_exp_syn;
wire o_LDPC_DEC_EXPSYND_78_exp_syn;
wire o_LDPC_DEC_EXPSYND_79_exp_syn;
wire o_LDPC_DEC_EXPSYND_80_exp_syn;
wire o_LDPC_DEC_EXPSYND_81_exp_syn;
wire o_LDPC_DEC_EXPSYND_82_exp_syn;
wire o_LDPC_DEC_EXPSYND_83_exp_syn;
wire o_LDPC_DEC_EXPSYND_84_exp_syn;
wire o_LDPC_DEC_EXPSYND_85_exp_syn;
wire o_LDPC_DEC_EXPSYND_86_exp_syn;
wire o_LDPC_DEC_EXPSYND_87_exp_syn;
wire o_LDPC_DEC_EXPSYND_88_exp_syn;
wire o_LDPC_DEC_EXPSYND_89_exp_syn;
wire o_LDPC_DEC_EXPSYND_90_exp_syn;
wire o_LDPC_DEC_EXPSYND_91_exp_syn;
wire o_LDPC_DEC_EXPSYND_92_exp_syn;
wire o_LDPC_DEC_EXPSYND_93_exp_syn;
wire o_LDPC_DEC_EXPSYND_94_exp_syn;
wire o_LDPC_DEC_EXPSYND_95_exp_syn;
wire o_LDPC_DEC_EXPSYND_96_exp_syn;
wire o_LDPC_DEC_EXPSYND_97_exp_syn;
wire o_LDPC_DEC_EXPSYND_98_exp_syn;
wire o_LDPC_DEC_EXPSYND_99_exp_syn;
wire o_LDPC_DEC_EXPSYND_100_exp_syn;
wire o_LDPC_DEC_EXPSYND_101_exp_syn;
wire o_LDPC_DEC_EXPSYND_102_exp_syn;
wire o_LDPC_DEC_EXPSYND_103_exp_syn;
wire o_LDPC_DEC_EXPSYND_104_exp_syn;
wire o_LDPC_DEC_EXPSYND_105_exp_syn;
wire o_LDPC_DEC_EXPSYND_106_exp_syn;
wire o_LDPC_DEC_EXPSYND_107_exp_syn;
wire o_LDPC_DEC_EXPSYND_108_exp_syn;
wire o_LDPC_DEC_EXPSYND_109_exp_syn;
wire o_LDPC_DEC_EXPSYND_110_exp_syn;
wire o_LDPC_DEC_EXPSYND_111_exp_syn;
wire o_LDPC_DEC_EXPSYND_112_exp_syn;
wire o_LDPC_DEC_EXPSYND_113_exp_syn;
wire o_LDPC_DEC_EXPSYND_114_exp_syn;
wire o_LDPC_DEC_EXPSYND_115_exp_syn;
wire o_LDPC_DEC_EXPSYND_116_exp_syn;
wire o_LDPC_DEC_EXPSYND_117_exp_syn;
wire o_LDPC_DEC_EXPSYND_118_exp_syn;
wire o_LDPC_DEC_EXPSYND_119_exp_syn;
wire o_LDPC_DEC_EXPSYND_120_exp_syn;
wire o_LDPC_DEC_EXPSYND_121_exp_syn;
wire o_LDPC_DEC_EXPSYND_122_exp_syn;
wire o_LDPC_DEC_EXPSYND_123_exp_syn;
wire o_LDPC_DEC_EXPSYND_124_exp_syn;
wire o_LDPC_DEC_EXPSYND_125_exp_syn;
wire o_LDPC_DEC_EXPSYND_126_exp_syn;
wire o_LDPC_DEC_EXPSYND_127_exp_syn;
wire o_LDPC_DEC_EXPSYND_128_exp_syn;
wire o_LDPC_DEC_EXPSYND_129_exp_syn;
wire o_LDPC_DEC_EXPSYND_130_exp_syn;
wire o_LDPC_DEC_EXPSYND_131_exp_syn;
wire o_LDPC_DEC_EXPSYND_132_exp_syn;
wire o_LDPC_DEC_EXPSYND_133_exp_syn;
wire o_LDPC_DEC_EXPSYND_134_exp_syn;
wire o_LDPC_DEC_EXPSYND_135_exp_syn;
wire o_LDPC_DEC_EXPSYND_136_exp_syn;
wire o_LDPC_DEC_EXPSYND_137_exp_syn;
wire o_LDPC_DEC_EXPSYND_138_exp_syn;
wire o_LDPC_DEC_EXPSYND_139_exp_syn;
wire o_LDPC_DEC_EXPSYND_140_exp_syn;
wire o_LDPC_DEC_EXPSYND_141_exp_syn;
wire o_LDPC_DEC_EXPSYND_142_exp_syn;
wire o_LDPC_DEC_EXPSYND_143_exp_syn;
wire o_LDPC_DEC_EXPSYND_144_exp_syn;
wire o_LDPC_DEC_EXPSYND_145_exp_syn;
wire o_LDPC_DEC_EXPSYND_146_exp_syn;
wire o_LDPC_DEC_EXPSYND_147_exp_syn;
wire o_LDPC_DEC_EXPSYND_148_exp_syn;
wire o_LDPC_DEC_EXPSYND_149_exp_syn;
wire o_LDPC_DEC_EXPSYND_150_exp_syn;
wire o_LDPC_DEC_EXPSYND_151_exp_syn;
wire o_LDPC_DEC_EXPSYND_152_exp_syn;
wire o_LDPC_DEC_EXPSYND_153_exp_syn;
wire o_LDPC_DEC_EXPSYND_154_exp_syn;
wire o_LDPC_DEC_EXPSYND_155_exp_syn;
wire o_LDPC_DEC_EXPSYND_156_exp_syn;
wire o_LDPC_DEC_EXPSYND_157_exp_syn;
wire o_LDPC_DEC_EXPSYND_158_exp_syn;
wire o_LDPC_DEC_EXPSYND_159_exp_syn;
wire o_LDPC_DEC_EXPSYND_160_exp_syn;
wire o_LDPC_DEC_EXPSYND_161_exp_syn;
wire o_LDPC_DEC_EXPSYND_162_exp_syn;
wire o_LDPC_DEC_EXPSYND_163_exp_syn;
wire o_LDPC_DEC_EXPSYND_164_exp_syn;
wire o_LDPC_DEC_EXPSYND_165_exp_syn;
wire o_LDPC_DEC_EXPSYND_166_exp_syn;
wire o_LDPC_DEC_EXPSYND_167_exp_syn;
wire [31:0] o_LDPC_DEC_PROBABILITY_perc_probability;
wire [31:0] o_LDPC_DEC_HAMDIST_LOOP_MAX_HamDist_loop_max;
wire [31:0] o_LDPC_DEC_HAMDIST_LOOP_PERCENTAGE_HamDist_loop_percentage;
wire [31:0] o_LDPC_DEC_HAMDIST_IIR1_HamDist_iir1;
wire [31:0] o_LDPC_DEC_HAMDIST_IIR2_NOT_USED_HamDist_iir2;
wire [31:0] o_LDPC_DEC_HAMDIST_IIR3_NOT_USED_HamDist_iir3;
wire i_LDPC_DEC_SYN_VALID_CWORD_DEC_NOT_USED_syn_valid_cword_dec;
wire o_LDPC_DEC_START_DEC_start_dec;
wire i_LDPC_DEC_CONVERGED_LOOPS_ENDED_converged_loops_ended;
wire i_LDPC_DEC_CONVERGED_PASS_FAIL_converged_pass_fail;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_0_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_1_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_2_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_3_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_4_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_5_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_6_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_7_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_8_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_9_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_10_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_11_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_12_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_13_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_14_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_15_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_16_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_17_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_18_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_19_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_20_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_21_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_22_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_23_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_24_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_25_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_26_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_27_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_28_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_29_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_30_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_31_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_32_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_33_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_34_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_35_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_36_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_37_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_38_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_39_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_40_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_41_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_42_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_43_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_44_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_45_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_46_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_47_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_48_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_49_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_50_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_51_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_52_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_53_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_54_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_55_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_56_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_57_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_58_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_59_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_60_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_61_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_62_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_63_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_64_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_65_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_66_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_67_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_68_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_69_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_70_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_71_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_72_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_73_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_74_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_75_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_76_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_77_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_78_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_79_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_80_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_81_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_82_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_83_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_84_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_85_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_86_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_87_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_88_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_89_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_90_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_91_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_92_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_93_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_94_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_95_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_96_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_97_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_98_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_99_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_100_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_101_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_102_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_103_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_104_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_105_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_106_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_107_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_108_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_109_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_110_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_111_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_112_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_113_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_114_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_115_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_116_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_117_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_118_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_119_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_120_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_121_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_122_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_123_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_124_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_125_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_126_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_127_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_128_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_129_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_130_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_131_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_132_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_133_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_134_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_135_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_136_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_137_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_138_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_139_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_140_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_141_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_142_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_143_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_144_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_145_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_146_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_147_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_148_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_149_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_150_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_151_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_152_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_153_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_154_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_155_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_156_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_157_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_158_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_159_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_160_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_161_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_162_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_163_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_164_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_165_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_166_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_167_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_168_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_169_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_170_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_171_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_172_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_173_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_174_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_175_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_176_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_177_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_178_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_179_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_180_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_181_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_182_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_183_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_184_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_185_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_186_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_187_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_188_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_189_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_190_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_191_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_192_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_193_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_194_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_195_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_196_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_197_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_198_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_199_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_200_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_201_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_202_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_203_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_204_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_205_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_206_final_cword;
wire i_LDPC_DEC_CODEWRD_OUT_BIT_207_final_cword;
wire o_LDPC_DEC_PASS_FAIL_pass_fail;
